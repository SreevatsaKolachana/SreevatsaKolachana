* PEX netlist file	Mon Apr 14 02:42:51 2025	Write_Driver
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 2
.subckt invx4 2 3 4 5 6 7 8
*.floating_nets 9 10 11 12
.ends invx4
.subckt sram_filler 2 3 4 5 6
.ends sram_filler
.subckt inv 2 3 4 5 6 8 9 10
*.floating_nets 7 11 12
MM1 3 5 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=395  $PIN_XY=420,380,390,395,360,380 $DEVICE_ID=1003
MM2 4 5 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=294  $PIN_XY=252,380,222,294,192,380 $DEVICE_ID=1003
.ends inv

* Hierarchy Level 1
.subckt buffer 2 3 4 5 6 7 8 9 10 11
XXACE67BBE10 2 3 5 4 7 9 10 11 inv $T=584 2 0 0 $X=584 $Y=2
XXACE67BBE11 2 3 4 6 8 9 10 11 inv $T=80 2 0 0 $X=80 $Y=2
.ends buffer
.subckt buffer_highdrive 2 3 4 5 6 7 8 9 10 11
MM1 2 5 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1568 $Y=393  $PIN_XY=1598,378,1568,393,1538,378 $DEVICE_ID=1003
MM2 4 5 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1400 $Y=393  $PIN_XY=1430,378,1400,393,1370,378 $DEVICE_ID=1003
MM3 2 5 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1232 $Y=313  $PIN_XY=1262,378,1232,313,1202,378 $DEVICE_ID=1003
MM4 4 5 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1064 $Y=313  $PIN_XY=1094,378,1064,313,1034,378 $DEVICE_ID=1003
MM5 2 6 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=728 $Y=393  $PIN_XY=758,378,728,393,698,378 $DEVICE_ID=1003
MM6 5 6 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=560 $Y=393  $PIN_XY=590,378,560,393,530,378 $DEVICE_ID=1003
MM7 2 6 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=392 $Y=292  $PIN_XY=422,378,392,292,362,378 $DEVICE_ID=1003
MM8 5 6 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=224 $Y=292  $PIN_XY=254,378,224,292,194,378 $DEVICE_ID=1003
XXACE67BBE12 3 2 5 6 9 10 11 invx4 $T=-22 -2 0 0 $X=2 $Y=-2
XXACE67BBE13 3 2 4 5 9 10 11 invx4 $T=818 -2 0 0 $X=842 $Y=-2
.ends buffer_highdrive

* Hierarchy Level 0

* Top of hierarchy  cell=Write_Driver
.subckt Write_Driver GND! VDD! DIN 5 6 WBDATA WDATA
MM1 GND! 16 WDATA nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2386 $Y=831  $PIN_XY=2416,936,2386,831,2356,936 $DEVICE_ID=1001
MM2 WDATA 16 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2218 $Y=831  $PIN_XY=2248,936,2218,831,2188,936 $DEVICE_ID=1001
MM3 GND! 6 WBDATA nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1546 $Y=1314  $PIN_XY=1576,1230,1546,1314,1516,1230 $DEVICE_ID=1001
MM4 GND! 5 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1546 $Y=852  $PIN_XY=1576,936,1546,852,1516,936 $DEVICE_ID=1001
MM5 WBDATA 6 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1378 $Y=1314  $PIN_XY=1408,1230,1378,1314,1348,1230 $DEVICE_ID=1001
MM6 16 5 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1378 $Y=852  $PIN_XY=1408,936,1378,852,1348,936 $DEVICE_ID=1001
MM7 6 9 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=874 $Y=1314  $PIN_XY=904,1230,874,1314,844,1230 $DEVICE_ID=1001
MM8 5 10 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=874 $Y=852  $PIN_XY=904,936,874,852,844,936 $DEVICE_ID=1001
MM9 9 DIN GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=370 $Y=1314  $PIN_XY=400,1230,370,1314,340,1230 $DEVICE_ID=1001
MM10 10 DIN GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=370 $Y=852  $PIN_XY=400,936,370,852,340,936 $DEVICE_ID=1001
MM11 VDD! 6 WBDATA pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1882 $Y=1415  $PIN_XY=1912,1400,1882,1415,1852,1400 $DEVICE_ID=1003
MM12 WBDATA 6 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1714 $Y=1415  $PIN_XY=1744,1400,1714,1415,1684,1400 $DEVICE_ID=1003
MM13 VDD! 6 WBDATA pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1546 $Y=1314  $PIN_XY=1576,1400,1546,1314,1516,1400 $DEVICE_ID=1003
MM14 WBDATA 6 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1378 $Y=1314  $PIN_XY=1408,1400,1378,1314,1348,1400 $DEVICE_ID=1003
XXACE67BBE1 GND! VDD! WBDATA 6 11 12 14 invx4 $T=1132 1020 0 0 $X=1156 $Y=1020
XXACE67BBE2 GND! VDD! 11 13 15 sram_filler $T=3284 1146 0 180 $X=2836 $Y=556
XXACE67BBE3 GND! VDD! 11 12 14 sram_filler $T=3284 1020 1 180 $X=2836 $Y=1020
XXACE67BBE4 GND! VDD! 11 12 14 sram_filler $T=2948 1020 1 180 $X=2500 $Y=1020
XXACE67BBE5 GND! VDD! 11 12 14 sram_filler $T=2328 1020 0 0 $X=2332 $Y=1020
XXACE67BBE6 GND! VDD! 11 12 14 sram_filler $T=1992 1020 0 0 $X=1996 $Y=1020
XXACE67BBE7 GND! VDD! 10 5 DIN 9 DIN 11 13 15 buffer $T=68 1148 1 0 $X=148 $Y=556
XXACE67BBE8 GND! VDD! 9 6 DIN 10 DIN 11 12 14 buffer $T=68 1018 0 0 $X=148 $Y=1020
XXACE67BBE9 VDD! GND! WDATA 16 5 6 6 11 13 15 buffer_highdrive $T=1154 1144 1 0 $X=1156 $Y=556
.ends Write_Driver
