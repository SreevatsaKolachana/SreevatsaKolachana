* PEX netlist file	Wed Apr 16 23:57:56 2025	sram_6t
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 0

* Top of hierarchy  cell=sram_6t
.subckt sram_6t 2 3 4 5 6 7 8 9 10 11
*.floating_nets 12 13 14 15 16 17 18 _GENERATED_19
MM1 4 6 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=366 $Y=756  $PIN_XY=396,840,366,756,336,840 $DEVICE_ID=1001
MM2 8 9 6 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=366 $Y=207  $PIN_XY=396,210,366,207,336,210 $DEVICE_ID=1001
MM3 7 9 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=198 $Y=843  $PIN_XY=228,840,198,843,168,840 $DEVICE_ID=1001
MM4 6 7 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=198 $Y=294  $PIN_XY=228,210,198,294,168,210 $DEVICE_ID=1001
MM5 3 6 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=366 $Y=756  $PIN_XY=396,670,366,756,336,670 $DEVICE_ID=1003
MM6 6 7 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=198 $Y=294  $PIN_XY=228,380,198,294,168,380 $DEVICE_ID=1003
.ends sram_6t
