* PEX netlist file	Mon Apr 14 01:32:34 2025	buffer_highdrive
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 1
.subckt invx4 2 3 4 5 6 7 8
*.floating_nets 9 10 11 12 13 14 15 16 17 18
MM1 2 5 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=414 $Y=294  $PIN_XY=444,210,414,294,384,210 $DEVICE_ID=1001
MM2 4 5 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=246 $Y=294  $PIN_XY=276,210,246,294,216,210 $DEVICE_ID=1001
MM3 3 5 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=750 $Y=395  $PIN_XY=780,380,750,395,720,380 $DEVICE_ID=1003
MM4 4 5 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=582 $Y=395  $PIN_XY=612,380,582,395,552,380 $DEVICE_ID=1003
MM5 3 5 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=414 $Y=294  $PIN_XY=444,380,414,294,384,380 $DEVICE_ID=1003
MM6 4 5 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=246 $Y=294  $PIN_XY=276,380,246,294,216,380 $DEVICE_ID=1003
.ends invx4

* Hierarchy Level 0

* Top of hierarchy  cell=buffer_highdrive
.subckt buffer_highdrive VDD! GND! 4 5
XX2533910A1 GND! VDD! 5 _GENERATED_9 6 7 8 invx4 $T=-22 -2 0 0 $X=2 $Y=-2
XX2533910A2 GND! VDD! 4 5 6 7 8 invx4 $T=818 -2 0 0 $X=842 $Y=-2
.ends buffer_highdrive
