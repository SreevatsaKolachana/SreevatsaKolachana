* PEX netlist file	Thu Apr 17 16:46:01 2025	static_row_decoder_3by8
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 2
.subckt nand 2 3 4 5 6 7 8 9 10 11 14
+	15
*.floating_nets 12 13
.ends nand
.subckt sram_filler 2 3 4 5 6 7
.ends sram_filler
.subckt nor 2 3 4 5 6 7 8 9 10 11 12
+	13
.ends nor
.subckt inv 2 3 4 5 6 8 9
*.floating_nets 7
.ends inv
.subckt invx4 2 3 4 5 6 7
.ends invx4

* Hierarchy Level 1
.subckt buffer_highdrive 2 3 4 5 6 7 8 9 10 11 12
XXF64012D8130 3 2 5 6 11 12 invx4 $T=-22 -2 0 0 $X=2 $Y=-2
XXF64012D8131 3 2 4 5 11 12 invx4 $T=818 -2 0 0 $X=842 $Y=-2
.ends buffer_highdrive

* Hierarchy Level 0

* Top of hierarchy  cell=static_row_decoder_3by8
.subckt static_row_decoder_3by8 VDD! GND! 4 5 6 7 8 9 10 11 12
+	A0 A1 15 16 WLREF A2 19 20 21 22 23
+	24 25 26 27 28 29 30 31 32 33 34
+	35 36
*.floating_nets 94 95 96 97 98 99 100 101 102 103
MM1 GND! 66 67 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=884  $PIN_XY=3760,800,3730,884,3700,800 $DEVICE_ID=1001
MM2 GND! 68 69 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-40  $PIN_XY=3760,-124,3730,-40,3700,-124 $DEVICE_ID=1001
MM3 GND! 61 62 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-964  $PIN_XY=3760,-1048,3730,-964,3700,-1048 $DEVICE_ID=1001
MM4 GND! 59 60 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-1888  $PIN_XY=3760,-1972,3730,-1888,3700,-1972 $DEVICE_ID=1001
MM5 GND! 55 56 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-2812  $PIN_XY=3760,-2896,3730,-2812,3700,-2896 $DEVICE_ID=1001
MM6 GND! 64 65 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-3736  $PIN_XY=3760,-3820,3730,-3736,3700,-3820 $DEVICE_ID=1001
MM7 GND! 57 58 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-4660  $PIN_XY=3760,-4744,3730,-4660,3700,-4744 $DEVICE_ID=1001
MM8 67 66 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=884  $PIN_XY=3592,800,3562,884,3532,800 $DEVICE_ID=1001
MM9 69 68 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-40  $PIN_XY=3592,-124,3562,-40,3532,-124 $DEVICE_ID=1001
MM10 62 61 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-964  $PIN_XY=3592,-1048,3562,-964,3532,-1048 $DEVICE_ID=1001
MM11 60 59 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-1888  $PIN_XY=3592,-1972,3562,-1888,3532,-1972 $DEVICE_ID=1001
MM12 56 55 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-2812  $PIN_XY=3592,-2896,3562,-2812,3532,-2896 $DEVICE_ID=1001
MM13 65 64 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-3736  $PIN_XY=3592,-3820,3562,-3736,3532,-3820 $DEVICE_ID=1001
MM14 58 57 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-4660  $PIN_XY=3592,-4744,3562,-4660,3532,-4744 $DEVICE_ID=1001
MM15 GND! 36 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=1346  $PIN_XY=2920,1430,2890,1346,2860,1430 $DEVICE_ID=1001
MM16 GND! 11 66 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=884  $PIN_XY=2920,800,2890,884,2860,800 $DEVICE_ID=1001
MM17 GND! 35 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=422  $PIN_XY=2920,506,2890,422,2860,506 $DEVICE_ID=1001
MM18 GND! 10 68 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-40  $PIN_XY=2920,-124,2890,-40,2860,-124 $DEVICE_ID=1001
MM19 GND! 34 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-502  $PIN_XY=2920,-418,2890,-502,2860,-418 $DEVICE_ID=1001
MM20 GND! 9 61 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-964  $PIN_XY=2920,-1048,2890,-964,2860,-1048 $DEVICE_ID=1001
MM21 GND! 33 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-1426  $PIN_XY=2920,-1342,2890,-1426,2860,-1342 $DEVICE_ID=1001
MM22 GND! 8 59 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-1888  $PIN_XY=2920,-1972,2890,-1888,2860,-1972 $DEVICE_ID=1001
MM23 GND! 27 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-2350  $PIN_XY=2920,-2266,2890,-2350,2860,-2266 $DEVICE_ID=1001
MM24 GND! 7 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-2812  $PIN_XY=2920,-2896,2890,-2812,2860,-2896 $DEVICE_ID=1001
MM25 GND! 26 6 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-3274  $PIN_XY=2920,-3190,2890,-3274,2860,-3190 $DEVICE_ID=1001
MM26 GND! 6 64 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-3736  $PIN_XY=2920,-3820,2890,-3736,2860,-3820 $DEVICE_ID=1001
MM27 GND! 25 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-4198  $PIN_XY=2920,-4114,2890,-4198,2860,-4114 $DEVICE_ID=1001
MM28 11 32 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=1346  $PIN_XY=2752,1430,2722,1346,2692,1430 $DEVICE_ID=1001
MM29 66 11 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=884  $PIN_XY=2752,800,2722,884,2692,800 $DEVICE_ID=1001
MM30 10 31 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=422  $PIN_XY=2752,506,2722,422,2692,506 $DEVICE_ID=1001
MM31 68 10 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-40  $PIN_XY=2752,-124,2722,-40,2692,-124 $DEVICE_ID=1001
MM32 9 30 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-502  $PIN_XY=2752,-418,2722,-502,2692,-418 $DEVICE_ID=1001
MM33 61 9 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-964  $PIN_XY=2752,-1048,2722,-964,2692,-1048 $DEVICE_ID=1001
MM34 8 29 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-1426  $PIN_XY=2752,-1342,2722,-1426,2692,-1342 $DEVICE_ID=1001
MM35 59 8 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-1888  $PIN_XY=2752,-1972,2722,-1888,2692,-1972 $DEVICE_ID=1001
MM36 7 23 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-2350  $PIN_XY=2752,-2266,2722,-2350,2692,-2266 $DEVICE_ID=1001
MM37 55 7 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-2812  $PIN_XY=2752,-2896,2722,-2812,2692,-2896 $DEVICE_ID=1001
MM38 6 22 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-3274  $PIN_XY=2752,-3190,2722,-3274,2692,-3190 $DEVICE_ID=1001
MM39 64 6 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-3736  $PIN_XY=2752,-3820,2722,-3736,2692,-3820 $DEVICE_ID=1001
MM40 5 21 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-4198  $PIN_XY=2752,-4114,2722,-4198,2692,-4114 $DEVICE_ID=1001
MM41 36 19 84 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=1346  $PIN_XY=2248,1430,2218,1346,2188,1430 $DEVICE_ID=1001
MM42 32 12 85 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=884  $PIN_XY=2248,800,2218,884,2188,800 $DEVICE_ID=1001
MM43 35 19 83 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=422  $PIN_XY=2248,506,2218,422,2188,506 $DEVICE_ID=1001
MM44 31 12 78 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-40  $PIN_XY=2248,-124,2218,-40,2188,-124 $DEVICE_ID=1001
MM45 34 A1 81 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-502  $PIN_XY=2248,-418,2218,-502,2188,-418 $DEVICE_ID=1001
MM46 30 12 82 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-964  $PIN_XY=2248,-1048,2218,-964,2188,-1048 $DEVICE_ID=1001
MM47 33 A1 80 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-1426  $PIN_XY=2248,-1342,2218,-1426,2188,-1342 $DEVICE_ID=1001
MM48 29 12 79 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-1888  $PIN_XY=2248,-1972,2218,-1888,2188,-1972 $DEVICE_ID=1001
MM49 27 19 71 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-2350  $PIN_XY=2248,-2266,2218,-2350,2188,-2266 $DEVICE_ID=1001
MM50 23 12 70 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-2812  $PIN_XY=2248,-2896,2218,-2812,2188,-2896 $DEVICE_ID=1001
MM51 26 19 72 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-3274  $PIN_XY=2248,-3190,2218,-3274,2188,-3190 $DEVICE_ID=1001
MM52 22 12 73 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-3736  $PIN_XY=2248,-3820,2218,-3736,2188,-3820 $DEVICE_ID=1001
MM53 25 A1 76 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-4198  $PIN_XY=2248,-4114,2218,-4198,2188,-4114 $DEVICE_ID=1001
MM54 84 15 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=1346  $PIN_XY=2080,1430,2050,1346,2020,1430 $DEVICE_ID=1001
MM55 85 28 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=884  $PIN_XY=2080,800,2050,884,2020,800 $DEVICE_ID=1001
MM56 83 A0 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=422  $PIN_XY=2080,506,2050,422,2020,506 $DEVICE_ID=1001
MM57 78 28 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-40  $PIN_XY=2080,-124,2050,-40,2020,-124 $DEVICE_ID=1001
MM58 81 15 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-502  $PIN_XY=2080,-418,2050,-502,2020,-418 $DEVICE_ID=1001
MM59 82 28 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-964  $PIN_XY=2080,-1048,2050,-964,2020,-1048 $DEVICE_ID=1001
MM60 80 A0 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-1426  $PIN_XY=2080,-1342,2050,-1426,2020,-1342 $DEVICE_ID=1001
MM61 79 28 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-1888  $PIN_XY=2080,-1972,2050,-1888,2020,-1972 $DEVICE_ID=1001
MM62 71 15 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-2350  $PIN_XY=2080,-2266,2050,-2350,2020,-2266 $DEVICE_ID=1001
MM63 70 A2 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-2812  $PIN_XY=2080,-2896,2050,-2812,2020,-2896 $DEVICE_ID=1001
MM64 72 A2 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-3274  $PIN_XY=2080,-3190,2050,-3274,2020,-3190 $DEVICE_ID=1001
MM65 73 A0 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-3736  $PIN_XY=2080,-3820,2050,-3736,2020,-3820 $DEVICE_ID=1001
MM66 76 15 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-4198  $PIN_XY=2080,-4114,2050,-4198,2020,-4114 $DEVICE_ID=1001
MM67 15 A0 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1546 $Y=1346  $PIN_XY=1576,1430,1546,1346,1516,1430 $DEVICE_ID=1001
MM68 19 A1 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1546 $Y=884  $PIN_XY=1576,800,1546,884,1516,800 $DEVICE_ID=1001
MM69 28 A2 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1546 $Y=443  $PIN_XY=1576,506,1546,443,1516,506 $DEVICE_ID=1001
MM70 GND! 37 63 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-5605  $PIN_XY=3760,-5668,3730,-5605,3700,-5668 $DEVICE_ID=1001
MM71 63 37 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-5605  $PIN_XY=3592,-5668,3562,-5605,3532,-5668 $DEVICE_ID=1001
MM72 GND! 5 57 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-4660  $PIN_XY=2920,-4744,2890,-4660,2860,-4744 $DEVICE_ID=1001
MM73 GND! 24 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-5122  $PIN_XY=2920,-5038,2890,-5122,2860,-5038 $DEVICE_ID=1001
MM74 GND! 4 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-5584  $PIN_XY=2920,-5668,2890,-5584,2860,-5668 $DEVICE_ID=1001
MM75 57 5 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-4660  $PIN_XY=2752,-4744,2722,-4660,2692,-4744 $DEVICE_ID=1001
MM76 4 20 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-5122  $PIN_XY=2752,-5038,2722,-5122,2692,-5038 $DEVICE_ID=1001
MM77 37 4 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-5584  $PIN_XY=2752,-5668,2722,-5584,2692,-5668 $DEVICE_ID=1001
MM78 21 12 75 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-4660  $PIN_XY=2248,-4744,2218,-4660,2188,-4744 $DEVICE_ID=1001
MM79 24 A1 77 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-5122  $PIN_XY=2248,-5038,2218,-5122,2188,-5038 $DEVICE_ID=1001
MM80 20 12 74 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-5584  $PIN_XY=2248,-5668,2218,-5584,2188,-5668 $DEVICE_ID=1001
MM81 75 A2 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-4660  $PIN_XY=2080,-4744,2050,-4660,2020,-4744 $DEVICE_ID=1001
MM82 77 A2 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-5122  $PIN_XY=2080,-5038,2050,-5122,2020,-5038 $DEVICE_ID=1001
MM83 74 A0 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-5584  $PIN_XY=2080,-5668,2050,-5584,2020,-5668 $DEVICE_ID=1001
MM84 GND! WLREF 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1042 $Y=-4681  $PIN_XY=1072,-4744,1042,-4681,1012,-4744 $DEVICE_ID=1001
MM85 GND! 16 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1042 $Y=-5101  $PIN_XY=1072,-5038,1042,-5101,1012,-5038 $DEVICE_ID=1001
MM86 16 WLREF GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=874 $Y=-4681  $PIN_XY=904,-4744,874,-4681,844,-4744 $DEVICE_ID=1001
MM87 12 16 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=874 $Y=-5101  $PIN_XY=904,-5038,874,-5101,844,-5038 $DEVICE_ID=1001
MM88 VDD! 66 67 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=964  $PIN_XY=4096,970,4066,964,4036,970 $DEVICE_ID=1003
MM89 VDD! 68 69 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=40  $PIN_XY=4096,46,4066,40,4036,46 $DEVICE_ID=1003
MM90 VDD! 61 62 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-884  $PIN_XY=4096,-878,4066,-884,4036,-878 $DEVICE_ID=1003
MM91 VDD! 59 60 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-1808  $PIN_XY=4096,-1802,4066,-1808,4036,-1802 $DEVICE_ID=1003
MM92 VDD! 55 56 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-2732  $PIN_XY=4096,-2726,4066,-2732,4036,-2726 $DEVICE_ID=1003
MM93 VDD! 64 65 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-3656  $PIN_XY=4096,-3650,4066,-3656,4036,-3650 $DEVICE_ID=1003
MM94 VDD! 57 58 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-4580  $PIN_XY=4096,-4574,4066,-4580,4036,-4574 $DEVICE_ID=1003
MM95 67 66 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=964  $PIN_XY=3928,970,3898,964,3868,970 $DEVICE_ID=1003
MM96 69 68 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=40  $PIN_XY=3928,46,3898,40,3868,46 $DEVICE_ID=1003
MM97 62 61 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-884  $PIN_XY=3928,-878,3898,-884,3868,-878 $DEVICE_ID=1003
MM98 60 59 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-1808  $PIN_XY=3928,-1802,3898,-1808,3868,-1802 $DEVICE_ID=1003
MM99 56 55 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-2732  $PIN_XY=3928,-2726,3898,-2732,3868,-2726 $DEVICE_ID=1003
MM100 65 64 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-3656  $PIN_XY=3928,-3650,3898,-3656,3868,-3650 $DEVICE_ID=1003
MM101 58 57 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-4580  $PIN_XY=3928,-4574,3898,-4580,3868,-4574 $DEVICE_ID=1003
MM102 VDD! 66 67 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=884  $PIN_XY=3760,970,3730,884,3700,970 $DEVICE_ID=1003
MM103 VDD! 68 69 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-40  $PIN_XY=3760,46,3730,-40,3700,46 $DEVICE_ID=1003
MM104 VDD! 61 62 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-964  $PIN_XY=3760,-878,3730,-964,3700,-878 $DEVICE_ID=1003
MM105 VDD! 59 60 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-1888  $PIN_XY=3760,-1802,3730,-1888,3700,-1802 $DEVICE_ID=1003
MM106 VDD! 55 56 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-2812  $PIN_XY=3760,-2726,3730,-2812,3700,-2726 $DEVICE_ID=1003
MM107 VDD! 64 65 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-3736  $PIN_XY=3760,-3650,3730,-3736,3700,-3650 $DEVICE_ID=1003
MM108 VDD! 57 58 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-4660  $PIN_XY=3760,-4574,3730,-4660,3700,-4574 $DEVICE_ID=1003
MM109 67 66 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=884  $PIN_XY=3592,970,3562,884,3532,970 $DEVICE_ID=1003
MM110 69 68 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-40  $PIN_XY=3592,46,3562,-40,3532,46 $DEVICE_ID=1003
MM111 62 61 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-964  $PIN_XY=3592,-878,3562,-964,3532,-878 $DEVICE_ID=1003
MM112 60 59 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-1888  $PIN_XY=3592,-1802,3562,-1888,3532,-1802 $DEVICE_ID=1003
MM113 56 55 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-2812  $PIN_XY=3592,-2726,3562,-2812,3532,-2726 $DEVICE_ID=1003
MM114 65 64 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-3736  $PIN_XY=3592,-3650,3562,-3736,3532,-3650 $DEVICE_ID=1003
MM115 58 57 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-4660  $PIN_XY=3592,-4574,3562,-4660,3532,-4574 $DEVICE_ID=1003
MM116 VDD! 11 66 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=964  $PIN_XY=3256,970,3226,964,3196,970 $DEVICE_ID=1003
MM117 VDD! 10 68 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=40  $PIN_XY=3256,46,3226,40,3196,46 $DEVICE_ID=1003
MM118 VDD! 9 61 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-884  $PIN_XY=3256,-878,3226,-884,3196,-878 $DEVICE_ID=1003
MM119 VDD! 8 59 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-1808  $PIN_XY=3256,-1802,3226,-1808,3196,-1802 $DEVICE_ID=1003
MM120 VDD! 7 55 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-2732  $PIN_XY=3256,-2726,3226,-2732,3196,-2726 $DEVICE_ID=1003
MM121 VDD! 6 64 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-3656  $PIN_XY=3256,-3650,3226,-3656,3196,-3650 $DEVICE_ID=1003
MM122 VDD! 5 57 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-4580  $PIN_XY=3256,-4574,3226,-4580,3196,-4574 $DEVICE_ID=1003
MM123 66 11 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=964  $PIN_XY=3088,970,3058,964,3028,970 $DEVICE_ID=1003
MM124 68 10 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=40  $PIN_XY=3088,46,3058,40,3028,46 $DEVICE_ID=1003
MM125 61 9 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-884  $PIN_XY=3088,-878,3058,-884,3028,-878 $DEVICE_ID=1003
MM126 59 8 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-1808  $PIN_XY=3088,-1802,3058,-1808,3028,-1802 $DEVICE_ID=1003
MM127 55 7 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-2732  $PIN_XY=3088,-2726,3058,-2732,3028,-2726 $DEVICE_ID=1003
MM128 64 6 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-3656  $PIN_XY=3088,-3650,3058,-3656,3028,-3650 $DEVICE_ID=1003
MM129 57 5 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-4580  $PIN_XY=3088,-4574,3058,-4580,3028,-4574 $DEVICE_ID=1003
MM130 11 36 92 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=1346  $PIN_XY=2920,1260,2890,1346,2860,1260 $DEVICE_ID=1003
MM131 VDD! 11 66 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=884  $PIN_XY=2920,970,2890,884,2860,970 $DEVICE_ID=1003
MM132 10 35 93 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=422  $PIN_XY=2920,336,2890,422,2860,336 $DEVICE_ID=1003
MM133 VDD! 10 68 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-40  $PIN_XY=2920,46,2890,-40,2860,46 $DEVICE_ID=1003
MM134 9 34 91 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-502  $PIN_XY=2920,-588,2890,-502,2860,-588 $DEVICE_ID=1003
MM135 VDD! 9 61 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-964  $PIN_XY=2920,-878,2890,-964,2860,-878 $DEVICE_ID=1003
MM136 8 33 90 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-1426  $PIN_XY=2920,-1512,2890,-1426,2860,-1512 $DEVICE_ID=1003
MM137 VDD! 8 59 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-1888  $PIN_XY=2920,-1802,2890,-1888,2860,-1802 $DEVICE_ID=1003
MM138 7 27 87 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-2350  $PIN_XY=2920,-2436,2890,-2350,2860,-2436 $DEVICE_ID=1003
MM139 VDD! 7 55 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-2812  $PIN_XY=2920,-2726,2890,-2812,2860,-2726 $DEVICE_ID=1003
MM140 6 26 88 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-3274  $PIN_XY=2920,-3360,2890,-3274,2860,-3360 $DEVICE_ID=1003
MM141 VDD! 6 64 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-3736  $PIN_XY=2920,-3650,2890,-3736,2860,-3650 $DEVICE_ID=1003
MM142 5 25 86 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-4198  $PIN_XY=2920,-4284,2890,-4198,2860,-4284 $DEVICE_ID=1003
MM143 92 32 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=1346  $PIN_XY=2752,1260,2722,1346,2692,1260 $DEVICE_ID=1003
MM144 66 11 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=884  $PIN_XY=2752,970,2722,884,2692,970 $DEVICE_ID=1003
MM145 93 31 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=422  $PIN_XY=2752,336,2722,422,2692,336 $DEVICE_ID=1003
MM146 68 10 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-40  $PIN_XY=2752,46,2722,-40,2692,46 $DEVICE_ID=1003
MM147 91 30 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-502  $PIN_XY=2752,-588,2722,-502,2692,-588 $DEVICE_ID=1003
MM148 61 9 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-964  $PIN_XY=2752,-878,2722,-964,2692,-878 $DEVICE_ID=1003
MM149 90 29 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-1426  $PIN_XY=2752,-1512,2722,-1426,2692,-1512 $DEVICE_ID=1003
MM150 59 8 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-1888  $PIN_XY=2752,-1802,2722,-1888,2692,-1802 $DEVICE_ID=1003
MM151 87 23 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-2350  $PIN_XY=2752,-2436,2722,-2350,2692,-2436 $DEVICE_ID=1003
MM152 55 7 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-2812  $PIN_XY=2752,-2726,2722,-2812,2692,-2726 $DEVICE_ID=1003
MM153 88 22 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-3274  $PIN_XY=2752,-3360,2722,-3274,2692,-3360 $DEVICE_ID=1003
MM154 64 6 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-3736  $PIN_XY=2752,-3650,2722,-3736,2692,-3650 $DEVICE_ID=1003
MM155 86 21 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-4198  $PIN_XY=2752,-4284,2722,-4198,2692,-4284 $DEVICE_ID=1003
MM156 VDD! 19 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=1346  $PIN_XY=2248,1260,2218,1346,2188,1260 $DEVICE_ID=1003
MM157 VDD! 12 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=884  $PIN_XY=2248,970,2218,884,2188,970 $DEVICE_ID=1003
MM158 VDD! 19 35 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=422  $PIN_XY=2248,336,2218,422,2188,336 $DEVICE_ID=1003
MM159 VDD! 12 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-40  $PIN_XY=2248,46,2218,-40,2188,46 $DEVICE_ID=1003
MM160 VDD! A1 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-502  $PIN_XY=2248,-588,2218,-502,2188,-588 $DEVICE_ID=1003
MM161 VDD! 12 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-964  $PIN_XY=2248,-878,2218,-964,2188,-878 $DEVICE_ID=1003
MM162 VDD! A1 33 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-1426  $PIN_XY=2248,-1512,2218,-1426,2188,-1512 $DEVICE_ID=1003
MM163 VDD! 12 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-1888  $PIN_XY=2248,-1802,2218,-1888,2188,-1802 $DEVICE_ID=1003
MM164 VDD! 19 27 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-2350  $PIN_XY=2248,-2436,2218,-2350,2188,-2436 $DEVICE_ID=1003
MM165 VDD! 12 23 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-2812  $PIN_XY=2248,-2726,2218,-2812,2188,-2726 $DEVICE_ID=1003
MM166 VDD! 19 26 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-3274  $PIN_XY=2248,-3360,2218,-3274,2188,-3360 $DEVICE_ID=1003
MM167 VDD! 12 22 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-3736  $PIN_XY=2248,-3650,2218,-3736,2188,-3650 $DEVICE_ID=1003
MM168 VDD! A1 25 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-4198  $PIN_XY=2248,-4284,2218,-4198,2188,-4284 $DEVICE_ID=1003
MM169 36 15 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=1346  $PIN_XY=2080,1260,2050,1346,2020,1260 $DEVICE_ID=1003
MM170 32 28 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=884  $PIN_XY=2080,970,2050,884,2020,970 $DEVICE_ID=1003
MM171 35 A0 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=422  $PIN_XY=2080,336,2050,422,2020,336 $DEVICE_ID=1003
MM172 31 28 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-40  $PIN_XY=2080,46,2050,-40,2020,46 $DEVICE_ID=1003
MM173 34 15 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-502  $PIN_XY=2080,-588,2050,-502,2020,-588 $DEVICE_ID=1003
MM174 30 28 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-964  $PIN_XY=2080,-878,2050,-964,2020,-878 $DEVICE_ID=1003
MM175 33 A0 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-1426  $PIN_XY=2080,-1512,2050,-1426,2020,-1512 $DEVICE_ID=1003
MM176 29 28 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-1888  $PIN_XY=2080,-1802,2050,-1888,2020,-1802 $DEVICE_ID=1003
MM177 27 15 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-2350  $PIN_XY=2080,-2436,2050,-2350,2020,-2436 $DEVICE_ID=1003
MM178 23 A2 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-2812  $PIN_XY=2080,-2726,2050,-2812,2020,-2726 $DEVICE_ID=1003
MM179 26 A2 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-3274  $PIN_XY=2080,-3360,2050,-3274,2020,-3360 $DEVICE_ID=1003
MM180 22 A0 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-3736  $PIN_XY=2080,-3650,2050,-3736,2020,-3650 $DEVICE_ID=1003
MM181 25 15 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-4198  $PIN_XY=2080,-4284,2050,-4198,2020,-4284 $DEVICE_ID=1003
MM182 VDD! A0 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1714 $Y=1245  $PIN_XY=1744,1260,1714,1245,1684,1260 $DEVICE_ID=1003
MM183 VDD! A1 19 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1714 $Y=985  $PIN_XY=1744,970,1714,985,1684,970 $DEVICE_ID=1003
MM184 VDD! A2 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1714 $Y=342  $PIN_XY=1744,336,1714,342,1684,336 $DEVICE_ID=1003
MM185 15 A0 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1546 $Y=1346  $PIN_XY=1576,1260,1546,1346,1516,1260 $DEVICE_ID=1003
MM186 19 A1 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1546 $Y=884  $PIN_XY=1576,970,1546,884,1516,970 $DEVICE_ID=1003
MM187 28 A2 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1546 $Y=443  $PIN_XY=1576,336,1546,443,1516,336 $DEVICE_ID=1003
MM188 VDD! WLREF 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1378 $Y=-4580  $PIN_XY=1408,-4574,1378,-4580,1348,-4574 $DEVICE_ID=1003
MM189 16 WLREF VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1210 $Y=-4580  $PIN_XY=1240,-4574,1210,-4580,1180,-4574 $DEVICE_ID=1003
MM190 VDD! 37 63 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-5504  $PIN_XY=4096,-5498,4066,-5504,4036,-5498 $DEVICE_ID=1003
MM191 63 37 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-5504  $PIN_XY=3928,-5498,3898,-5504,3868,-5498 $DEVICE_ID=1003
MM192 VDD! 37 63 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-5605  $PIN_XY=3760,-5498,3730,-5605,3700,-5498 $DEVICE_ID=1003
MM193 63 37 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-5605  $PIN_XY=3592,-5498,3562,-5605,3532,-5498 $DEVICE_ID=1003
MM194 VDD! 4 37 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-5504  $PIN_XY=3256,-5498,3226,-5504,3196,-5498 $DEVICE_ID=1003
MM195 37 4 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-5504  $PIN_XY=3088,-5498,3058,-5504,3028,-5498 $DEVICE_ID=1003
MM196 VDD! 5 57 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-4660  $PIN_XY=2920,-4574,2890,-4660,2860,-4574 $DEVICE_ID=1003
MM197 4 24 89 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-5122  $PIN_XY=2920,-5208,2890,-5122,2860,-5208 $DEVICE_ID=1003
MM198 VDD! 4 37 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-5584  $PIN_XY=2920,-5498,2890,-5584,2860,-5498 $DEVICE_ID=1003
MM199 57 5 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-4660  $PIN_XY=2752,-4574,2722,-4660,2692,-4574 $DEVICE_ID=1003
MM200 89 20 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-5122  $PIN_XY=2752,-5208,2722,-5122,2692,-5208 $DEVICE_ID=1003
MM201 37 4 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-5584  $PIN_XY=2752,-5498,2722,-5584,2692,-5498 $DEVICE_ID=1003
MM202 VDD! 12 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-4660  $PIN_XY=2248,-4574,2218,-4660,2188,-4574 $DEVICE_ID=1003
MM203 VDD! A1 24 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-5122  $PIN_XY=2248,-5208,2218,-5122,2188,-5208 $DEVICE_ID=1003
MM204 VDD! 12 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-5584  $PIN_XY=2248,-5498,2218,-5584,2188,-5498 $DEVICE_ID=1003
MM205 21 A2 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-4660  $PIN_XY=2080,-4574,2050,-4660,2020,-4574 $DEVICE_ID=1003
MM206 24 A2 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-5122  $PIN_XY=2080,-5208,2050,-5122,2020,-5208 $DEVICE_ID=1003
MM207 20 A0 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-5584  $PIN_XY=2080,-5498,2050,-5584,2020,-5498 $DEVICE_ID=1003
MM208 VDD! 16 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1378 $Y=-5202  $PIN_XY=1408,-5208,1378,-5202,1348,-5208 $DEVICE_ID=1003
MM209 12 16 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1210 $Y=-5202  $PIN_XY=1240,-5208,1210,-5202,1180,-5208 $DEVICE_ID=1003
MM210 VDD! WLREF 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1042 $Y=-4681  $PIN_XY=1072,-4574,1042,-4681,1012,-4574 $DEVICE_ID=1003
MM211 VDD! 16 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1042 $Y=-5101  $PIN_XY=1072,-5208,1042,-5101,1012,-5208 $DEVICE_ID=1003
MM212 16 WLREF VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=874 $Y=-4681  $PIN_XY=904,-4574,874,-4681,844,-4574 $DEVICE_ID=1003
MM213 12 16 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=874 $Y=-5101  $PIN_XY=904,-5208,874,-5101,844,-5208 $DEVICE_ID=1003
XXF64012D81 VDD! GND! 56 55 7 22 23 26 27 40 50 buffer_highdrive $T=2498 -3104 0 0 $X=2500 $Y=-3106
XXF64012D82 VDD! GND! 58 57 5 20 21 24 25 39 48 buffer_highdrive $T=2498 -4952 0 0 $X=2500 $Y=-4954
XXF64012D83 VDD! GND! 60 59 8 23 29 27 33 43 51 buffer_highdrive $T=2498 -2180 0 0 $X=2500 $Y=-2182
XXF64012D84 VDD! GND! 62 61 9 29 30 33 34 42 53 buffer_highdrive $T=2498 -1256 0 0 $X=2500 $Y=-1258
XXF64012D85 VDD! GND! 63 37 4 106 20 107 24 38 47 buffer_highdrive $T=2498 -5876 0 0 $X=2500 $Y=-5878
XXF64012D86 VDD! GND! 65 64 6 21 22 25 26 41 49 buffer_highdrive $T=2498 -4028 0 0 $X=2500 $Y=-4030
XXF64012D87 VDD! GND! 67 66 11 31 32 35 36 45 54 buffer_highdrive $T=2498 592 0 0 $X=2500 $Y=590
XXF64012D88 VDD! GND! 69 68 10 30 31 34 35 46 52 buffer_highdrive $T=2498 -332 0 0 $X=2500 $Y=-334
XXF64012D89 GND! VDD! 12 16 39 47 invx4 $T=628 -4828 1 0 $X=652 $Y=-5418
XXF64012D810 GND! VDD! 16 WLREF 39 48 invx4 $T=628 -4954 0 0 $X=652 $Y=-4954
XXF64012D811 GND! VDD! _GENERATED_114 _GENERATED_113 42 53 sram_filler $T=4176 -1258 0 0 $X=4180 $Y=-1258
XXF64012D812 GND! VDD! _GENERATED_116 _GENERATED_115 40 49 sram_filler $T=4628 -2980 0 180 $X=4180 $Y=-3570
XXF64012D813 GND! VDD! _GENERATED_118 _GENERATED_117 40 50 sram_filler $T=4176 -3106 0 0 $X=4180 $Y=-3106
XXF64012D814 GND! VDD! _GENERATED_120 _GENERATED_119 43 50 sram_filler $T=4628 -2056 0 180 $X=4180 $Y=-2646
XXF64012D815 GND! VDD! _GENERATED_122 _GENERATED_121 43 51 sram_filler $T=4176 -2182 0 0 $X=4180 $Y=-2182
XXF64012D816 GND! VDD! _GENERATED_124 _GENERATED_123 42 51 sram_filler $T=4628 -1132 0 180 $X=4180 $Y=-1722
XXF64012D817 GND! VDD! _GENERATED_126 _GENERATED_125 41 49 sram_filler $T=4176 -4030 0 0 $X=4180 $Y=-4030
XXF64012D818 GND! VDD! _GENERATED_128 _GENERATED_127 41 48 sram_filler $T=4628 -3904 0 180 $X=4180 $Y=-4494
XXF64012D819 GND! VDD! _GENERATED_130 _GENERATED_129 39 48 sram_filler $T=4176 -4954 0 0 $X=4180 $Y=-4954
XXF64012D820 GND! VDD! _GENERATED_132 _GENERATED_131 39 47 sram_filler $T=4628 -4828 0 180 $X=4180 $Y=-5418
XXF64012D821 GND! VDD! _GENERATED_134 _GENERATED_133 38 47 sram_filler $T=4176 -5878 0 0 $X=4180 $Y=-5878
XXF64012D822 GND! VDD! _GENERATED_136 _GENERATED_135 46 53 sram_filler $T=4628 -208 0 180 $X=4180 $Y=-798
XXF64012D823 GND! VDD! _GENERATED_138 _GENERATED_137 46 52 sram_filler $T=4176 -334 0 0 $X=4180 $Y=-334
XXF64012D824 GND! VDD! _GENERATED_140 _GENERATED_139 45 52 sram_filler $T=4628 716 0 180 $X=4180 $Y=126
XXF64012D825 GND! VDD! _GENERATED_142 _GENERATED_141 45 54 sram_filler $T=4176 590 0 0 $X=4180 $Y=590
XXF64012D826 GND! VDD! _GENERATED_144 _GENERATED_143 44 54 sram_filler $T=4628 1640 0 180 $X=4180 $Y=1050
XXF64012D827 GND! VDD! _GENERATED_146 _GENERATED_145 44 54 sram_filler $T=1100 1640 0 180 $X=652 $Y=1050
XXF64012D828 GND! VDD! _GENERATED_148 _GENERATED_147 45 54 sram_filler $T=648 590 0 0 $X=652 $Y=590
XXF64012D829 GND! VDD! _GENERATED_150 _GENERATED_149 45 52 sram_filler $T=1100 716 0 180 $X=652 $Y=126
XXF64012D830 GND! VDD! _GENERATED_152 _GENERATED_151 45 52 sram_filler $T=1436 716 0 180 $X=988 $Y=126
XXF64012D831 GND! VDD! _GENERATED_154 _GENERATED_153 45 54 sram_filler $T=984 590 0 0 $X=988 $Y=590
XXF64012D832 GND! VDD! _GENERATED_156 _GENERATED_155 44 54 sram_filler $T=1436 1640 0 180 $X=988 $Y=1050
XXF64012D833 GND! VDD! _GENERATED_158 _GENERATED_157 38 47 sram_filler $T=648 -5878 0 0 $X=652 $Y=-5878
XXF64012D834 GND! VDD! _GENERATED_160 _GENERATED_159 38 47 sram_filler $T=984 -5878 0 0 $X=988 $Y=-5878
XXF64012D835 GND! VDD! _GENERATED_161 GND! 38 47 sram_filler $T=1320 -5878 0 0 $X=1324 $Y=-5878
XXF64012D836 GND! VDD! VDD! _GENERATED_162 38 47 sram_filler $T=1488 -5878 0 0 $X=1492 $Y=-5878
XXF64012D837 GND! VDD! _GENERATED_164 _GENERATED_163 46 52 sram_filler $T=648 -334 0 0 $X=652 $Y=-334
XXF64012D838 GND! VDD! _GENERATED_166 _GENERATED_165 46 52 sram_filler $T=984 -334 0 0 $X=988 $Y=-334
XXF64012D839 GND! VDD! _GENERATED_167 GND! 46 52 sram_filler $T=1320 -334 0 0 $X=1324 $Y=-334
XXF64012D840 GND! VDD! VDD! _GENERATED_168 46 52 sram_filler $T=1488 -334 0 0 $X=1492 $Y=-334
XXF64012D841 GND! VDD! _GENERATED_169 GND! 42 53 sram_filler $T=648 -1258 0 0 $X=652 $Y=-1258
XXF64012D842 GND! VDD! VDD! _GENERATED_170 42 53 sram_filler $T=816 -1258 0 0 $X=820 $Y=-1258
XXF64012D843 GND! VDD! _GENERATED_172 _GENERATED_171 42 53 sram_filler $T=1152 -1258 0 0 $X=1156 $Y=-1258
XXF64012D844 GND! VDD! _GENERATED_174 _GENERATED_173 42 53 sram_filler $T=1488 -1258 0 0 $X=1492 $Y=-1258
XXF64012D845 GND! VDD! VDD! _GENERATED_175 46 53 sram_filler $T=1100 -208 0 180 $X=652 $Y=-798
XXF64012D846 GND! VDD! _GENERATED_176 GND! 46 53 sram_filler $T=1268 -208 0 180 $X=820 $Y=-798
XXF64012D847 GND! VDD! _GENERATED_178 _GENERATED_177 46 53 sram_filler $T=1604 -208 0 180 $X=1156 $Y=-798
XXF64012D848 GND! VDD! _GENERATED_180 _GENERATED_179 46 53 sram_filler $T=1940 -208 0 180 $X=1492 $Y=-798
XXF64012D849 GND! VDD! _GENERATED_182 _GENERATED_181 42 51 sram_filler $T=1940 -1132 0 180 $X=1492 $Y=-1722
XXF64012D850 GND! VDD! _GENERATED_184 _GENERATED_183 42 51 sram_filler $T=1604 -1132 0 180 $X=1156 $Y=-1722
XXF64012D851 GND! VDD! _GENERATED_185 GND! 42 51 sram_filler $T=1268 -1132 0 180 $X=820 $Y=-1722
XXF64012D852 GND! VDD! VDD! _GENERATED_186 42 51 sram_filler $T=1100 -1132 0 180 $X=652 $Y=-1722
XXF64012D853 GND! VDD! _GENERATED_188 _GENERATED_187 43 51 sram_filler $T=1488 -2182 0 0 $X=1492 $Y=-2182
XXF64012D854 GND! VDD! _GENERATED_190 _GENERATED_189 43 51 sram_filler $T=1152 -2182 0 0 $X=1156 $Y=-2182
XXF64012D855 GND! VDD! VDD! _GENERATED_191 43 51 sram_filler $T=816 -2182 0 0 $X=820 $Y=-2182
XXF64012D856 GND! VDD! _GENERATED_192 GND! 43 51 sram_filler $T=648 -2182 0 0 $X=652 $Y=-2182
XXF64012D857 GND! VDD! VDD! _GENERATED_193 43 50 sram_filler $T=1100 -2056 0 180 $X=652 $Y=-2646
XXF64012D858 GND! VDD! _GENERATED_194 GND! 43 50 sram_filler $T=1268 -2056 0 180 $X=820 $Y=-2646
XXF64012D859 GND! VDD! _GENERATED_196 _GENERATED_195 43 50 sram_filler $T=1604 -2056 0 180 $X=1156 $Y=-2646
XXF64012D860 GND! VDD! _GENERATED_198 _GENERATED_197 43 50 sram_filler $T=1940 -2056 0 180 $X=1492 $Y=-2646
XXF64012D861 GND! VDD! _GENERATED_200 _GENERATED_199 40 50 sram_filler $T=648 -3106 0 0 $X=652 $Y=-3106
XXF64012D862 GND! VDD! _GENERATED_202 _GENERATED_201 40 50 sram_filler $T=984 -3106 0 0 $X=988 $Y=-3106
XXF64012D863 GND! VDD! _GENERATED_203 GND! 40 50 sram_filler $T=1320 -3106 0 0 $X=1324 $Y=-3106
XXF64012D864 GND! VDD! VDD! _GENERATED_204 40 50 sram_filler $T=1488 -3106 0 0 $X=1492 $Y=-3106
XXF64012D865 GND! VDD! _GENERATED_206 _GENERATED_205 40 49 sram_filler $T=1940 -2980 0 180 $X=1492 $Y=-3570
XXF64012D866 GND! VDD! _GENERATED_208 _GENERATED_207 40 49 sram_filler $T=1604 -2980 0 180 $X=1156 $Y=-3570
XXF64012D867 GND! VDD! _GENERATED_209 GND! 40 49 sram_filler $T=1268 -2980 0 180 $X=820 $Y=-3570
XXF64012D868 GND! VDD! VDD! _GENERATED_210 40 49 sram_filler $T=1100 -2980 0 180 $X=652 $Y=-3570
XXF64012D869 GND! VDD! VDD! _GENERATED_211 41 49 sram_filler $T=1488 -4030 0 0 $X=1492 $Y=-4030
XXF64012D870 GND! VDD! _GENERATED_212 GND! 41 49 sram_filler $T=1320 -4030 0 0 $X=1324 $Y=-4030
XXF64012D871 GND! VDD! _GENERATED_214 _GENERATED_213 41 49 sram_filler $T=984 -4030 0 0 $X=988 $Y=-4030
XXF64012D872 GND! VDD! _GENERATED_216 _GENERATED_215 41 49 sram_filler $T=648 -4030 0 0 $X=652 $Y=-4030
XXF64012D873 GND! VDD! VDD! _GENERATED_217 41 48 sram_filler $T=1100 -3904 0 180 $X=652 $Y=-4494
XXF64012D874 GND! VDD! _GENERATED_218 GND! 41 48 sram_filler $T=1268 -3904 0 180 $X=820 $Y=-4494
XXF64012D875 GND! VDD! _GENERATED_220 _GENERATED_219 41 48 sram_filler $T=1604 -3904 0 180 $X=1156 $Y=-4494
XXF64012D876 GND! VDD! _GENERATED_222 _GENERATED_221 41 48 sram_filler $T=1940 -3904 0 180 $X=1492 $Y=-4494
XXF64012D877 GND! VDD! _GENERATED_224 _GENERATED_223 43 50 sram_filler $T=3168 -2056 1 0 $X=3172 $Y=-2646
XXF64012D878 GND! VDD! _GENERATED_226 _GENERATED_225 43 50 sram_filler $T=3840 -2056 1 0 $X=3844 $Y=-2646
XXF64012D879 GND! VDD! _GENERATED_228 _GENERATED_227 43 50 sram_filler $T=3504 -2056 1 0 $X=3508 $Y=-2646
XXF64012D880 GND! VDD! _GENERATED_230 _GENERATED_229 40 49 sram_filler $T=3840 -2980 1 0 $X=3844 $Y=-3570
XXF64012D881 GND! VDD! _GENERATED_232 _GENERATED_231 40 49 sram_filler $T=3168 -2980 1 0 $X=3172 $Y=-3570
XXF64012D882 GND! VDD! _GENERATED_234 _GENERATED_233 40 49 sram_filler $T=3504 -2980 1 0 $X=3508 $Y=-3570
XXF64012D883 GND! VDD! _GENERATED_236 _GENERATED_235 41 48 sram_filler $T=3168 -3904 1 0 $X=3172 $Y=-4494
XXF64012D884 GND! VDD! _GENERATED_238 _GENERATED_237 41 48 sram_filler $T=3840 -3904 1 0 $X=3844 $Y=-4494
XXF64012D885 GND! VDD! _GENERATED_240 _GENERATED_239 41 48 sram_filler $T=3504 -3904 1 0 $X=3508 $Y=-4494
XXF64012D886 GND! VDD! _GENERATED_242 _GENERATED_241 39 47 sram_filler $T=3840 -4828 1 0 $X=3844 $Y=-5418
XXF64012D887 GND! VDD! _GENERATED_244 _GENERATED_243 39 47 sram_filler $T=3168 -4828 1 0 $X=3172 $Y=-5418
XXF64012D888 GND! VDD! _GENERATED_246 _GENERATED_245 39 47 sram_filler $T=3504 -4828 1 0 $X=3508 $Y=-5418
XXF64012D889 GND! VDD! _GENERATED_248 _GENERATED_247 42 51 sram_filler $T=3504 -1132 1 0 $X=3508 $Y=-1722
XXF64012D890 GND! VDD! _GENERATED_250 _GENERATED_249 42 51 sram_filler $T=3168 -1132 1 0 $X=3172 $Y=-1722
XXF64012D891 GND! VDD! _GENERATED_252 _GENERATED_251 42 51 sram_filler $T=3840 -1132 1 0 $X=3844 $Y=-1722
XXF64012D892 GND! VDD! _GENERATED_254 _GENERATED_253 46 53 sram_filler $T=3504 -208 1 0 $X=3508 $Y=-798
XXF64012D893 GND! VDD! _GENERATED_256 _GENERATED_255 46 53 sram_filler $T=3840 -208 1 0 $X=3844 $Y=-798
XXF64012D894 GND! VDD! _GENERATED_258 _GENERATED_257 46 53 sram_filler $T=3168 -208 1 0 $X=3172 $Y=-798
XXF64012D895 GND! VDD! _GENERATED_260 _GENERATED_259 45 52 sram_filler $T=3168 716 1 0 $X=3172 $Y=126
XXF64012D896 GND! VDD! _GENERATED_262 _GENERATED_261 45 52 sram_filler $T=3840 716 1 0 $X=3844 $Y=126
XXF64012D897 GND! VDD! _GENERATED_264 _GENERATED_263 44 54 sram_filler $T=3840 1640 1 0 $X=3844 $Y=1050
XXF64012D898 GND! VDD! _GENERATED_266 _GENERATED_265 44 54 sram_filler $T=3168 1640 1 0 $X=3172 $Y=1050
XXF64012D899 GND! VDD! _GENERATED_268 _GENERATED_267 44 54 sram_filler $T=3504 1640 1 0 $X=3508 $Y=1050
XXF64012D8100 GND! VDD! _GENERATED_270 _GENERATED_269 45 52 sram_filler $T=3504 716 1 0 $X=3508 $Y=126
XXF64012D8101 GND! VDD! _GENERATED_272 _GENERATED_271 39 47 sram_filler $T=1488 -4828 1 0 $X=1492 $Y=-5418
XXF64012D8102 GND! VDD! _GENERATED_274 _GENERATED_273 39 48 sram_filler $T=1488 -4954 0 0 $X=1492 $Y=-4954
XXF64012D8103 GND! VDD! 28 A2 A1 45 52 inv $T=1324 716 1 0 $X=1324 $Y=126
XXF64012D8104 GND! VDD! 15 A0 108 44 54 inv $T=1324 1640 1 0 $X=1324 $Y=1050
XXF64012D8105 GND! VDD! 19 A1 A2 45 54 inv $T=1324 590 0 0 $X=1324 $Y=590
XXF64012D8106 GND! VDD! 23 A2 12 A2 15 19 19 70 40 
+	50 nand $T=1410 -3334 0 0 $X=1827 $Y=-3106
XXF64012D8107 GND! VDD! 27 15 19 28 A2 12 12 71 43 
+	50 nand $T=1410 -1828 1 0 $X=1827 $Y=-2646
XXF64012D8108 GND! VDD! 26 A2 19 A2 A0 12 12 72 40 
+	49 nand $T=1410 -2752 1 0 $X=1827 $Y=-3570
XXF64012D8109 GND! VDD! 22 A0 12 15 A2 A1 19 73 41 
+	49 nand $T=1410 -4258 0 0 $X=1827 $Y=-4030
XXF64012D8110 GND! VDD! 20 A0 12 104 A2 105 A1 74 38 
+	47 nand $T=1410 -6106 0 0 $X=1827 $Y=-5878
XXF64012D8111 GND! VDD! 21 A2 12 A2 15 A1 A1 75 39 
+	48 nand $T=1410 -5182 0 0 $X=1827 $Y=-4954
XXF64012D8112 GND! VDD! 25 15 A1 A0 A2 12 12 76 41 
+	48 nand $T=1410 -3676 1 0 $X=1827 $Y=-4494
XXF64012D8113 GND! VDD! 24 A2 A1 A2 A0 12 12 77 39 
+	47 nand $T=1410 -4600 1 0 $X=1827 $Y=-5418
XXF64012D8114 GND! VDD! 31 28 12 15 A0 A1 19 78 46 
+	52 nand $T=1410 -562 0 0 $X=1827 $Y=-334
XXF64012D8115 GND! VDD! 29 28 12 15 A0 19 A1 79 43 
+	51 nand $T=1410 -2410 0 0 $X=1827 $Y=-2182
XXF64012D8116 GND! VDD! 33 A0 A1 28 28 12 12 80 42 
+	51 nand $T=1410 -904 1 0 $X=1827 $Y=-1722
XXF64012D8117 GND! VDD! 34 15 A1 28 28 12 12 81 46 
+	53 nand $T=1410 20 1 0 $X=1827 $Y=-798
XXF64012D8118 GND! VDD! 30 28 12 A0 15 A1 A1 82 42 
+	53 nand $T=1410 -1486 0 0 $X=1827 $Y=-1258
XXF64012D8119 GND! VDD! 35 A0 19 28 28 12 12 83 45 
+	52 nand $T=1410 944 1 0 $X=1827 $Y=126
XXF64012D8120 GND! VDD! 36 15 19 109 28 110 12 84 44 
+	54 nand $T=1410 1868 1 0 $X=1827 $Y=1050
XXF64012D8121 GND! VDD! 32 28 12 A0 15 19 19 85 45 
+	54 nand $T=1410 362 0 0 $X=1827 $Y=590
XXF64012D8122 GND! VDD! 5 21 25 6 5 6 5 86 41 
+	48 nor $T=1872 -3902 1 0 $X=2500 $Y=-4494
XXF64012D8123 GND! VDD! 7 23 27 8 7 8 7 87 43 
+	50 nor $T=1872 -2054 1 0 $X=2500 $Y=-2646
XXF64012D8124 GND! VDD! 6 22 26 7 6 7 6 88 40 
+	49 nor $T=1872 -2978 1 0 $X=2500 $Y=-3570
XXF64012D8125 GND! VDD! 4 20 24 5 4 5 4 89 39 
+	47 nor $T=1872 -4826 1 0 $X=2500 $Y=-5418
XXF64012D8126 GND! VDD! 8 29 33 9 8 9 8 90 42 
+	51 nor $T=1872 -1130 1 0 $X=2500 $Y=-1722
XXF64012D8127 GND! VDD! 9 30 34 10 9 10 9 91 46 
+	53 nor $T=1872 -206 1 0 $X=2500 $Y=-798
XXF64012D8128 GND! VDD! 11 32 36 111 11 112 11 92 44 
+	54 nor $T=1872 1642 1 0 $X=2500 $Y=1050
XXF64012D8129 GND! VDD! 10 31 35 11 10 11 10 93 45 
+	52 nor $T=1872 718 1 0 $X=2500 $Y=126
.ends static_row_decoder_3by8
