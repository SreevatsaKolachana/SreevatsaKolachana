* PEX netlist file	Fri Apr 18 03:45:02 2025	integration
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 3
.subckt sram_filler 2 3 4 5 6 7
.ends sram_filler
.subckt tspc_pos_ff 2 3 4 8 9 25 26 27
*.floating_nets 10 11 13 14 15 17 18 19 20 22 23
*+	24 28 29 30 31 32 33 34 35
MM1 4 7 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1176 $Y=294  $PIN_XY=1206,210,1176,294,1146,210 $DEVICE_ID=1001
MM2 2 6 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1008 $Y=294  $PIN_XY=1038,210,1008,294,978,210 $DEVICE_ID=1001
MM3 16 9 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=840 $Y=209  $PIN_XY=870,210,840,209,810,210 $DEVICE_ID=1001
MM4 6 9 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=504 $Y=209  $PIN_XY=534,210,504,209,474,210 $DEVICE_ID=1001
MM5 12 5 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=336 $Y=209  $PIN_XY=366,210,336,209,306,210 $DEVICE_ID=1001
MM6 2 8 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=168 $Y=209  $PIN_XY=198,210,168,209,138,210 $DEVICE_ID=1001
MM7 4 7 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1176 $Y=294  $PIN_XY=1206,380,1176,294,1146,380 $DEVICE_ID=1003
MM8 3 6 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1008 $Y=294  $PIN_XY=1038,380,1008,294,978,380 $DEVICE_ID=1003
MM9 5 9 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=504 $Y=649  $PIN_XY=534,670,504,649,474,670 $DEVICE_ID=1003
MM10 21 8 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=336 $Y=670  $PIN_XY=366,670,336,670,306,670 $DEVICE_ID=1003
MM11 3 9 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=168 $Y=670  $PIN_XY=198,670,168,670,138,670 $DEVICE_ID=1003
.ends tspc_pos_ff
.subckt nand 2 3 4 5 6 7 10 11
*.floating_nets 8 9
.ends nand
.subckt inv 2 3 4 5 7 8
*.floating_nets 6
.ends inv
.subckt 2to4_decoder_static_filler_17 2 3 4 5 6 7
.ends 2to4_decoder_static_filler_17
.subckt Filler 2 3 4 5 6 7 8 9
.ends Filler
.subckt precharge_logic 2 3 4 5 6 7 8 11 12
*.floating_nets 9 10
.ends precharge_logic
.subckt sram_6t 2 3 4 5 6 7 8 9 10 11 14
+	15 16
*.floating_nets 12 13 17 18
MM1 3 6 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=366 $Y=756  $PIN_XY=396,670,366,756,336,670 $DEVICE_ID=1003
.ends sram_6t
.subckt bitcell_precharge_filler 2 3 4 5 6 7
.ends bitcell_precharge_filler
.subckt nor 2 3 4 5 6 7 8 9
.ends nor
.subckt invx4 2 3 4 5 6 7
.ends invx4

* Hierarchy Level 2
.subckt 2to4_decoder_static 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16 17 18 19 20 21 22 25
+	27 29 30 32 34 36 38 39 40 41 42
+	43 44 45 46 79 80 81 82 83 84 85
+	86 87
*.floating_nets 47 48 49 50 51 52 53 54 55 56 57
*+	58 59 60 61 62 63 64 65 66 67 68
*+	69 70 71 72 73 74 75 76 77 78 96
*+	97 98 99 100 101 102 103
MM1 18 37 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2574 $Y=2243  $PIN_XY=2604,2226,2574,2243,2544,2226 $DEVICE_ID=1001
MM2 5 25 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=1197  $PIN_XY=2436,1302,2406,1197,2376,1302 $DEVICE_ID=1001
MM3 46 43 95 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=294  $PIN_XY=2436,378,2406,294,2376,378 $DEVICE_ID=1001
MM4 17 37 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2238 $Y=2244  $PIN_XY=2268,2226,2238,2244,2208,2226 $DEVICE_ID=1001
MM5 38 24 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2238 $Y=1680  $PIN_XY=2268,1596,2238,1680,2208,1596 $DEVICE_ID=1001
MM6 24 42 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=1218  $PIN_XY=2268,1302,2238,1218,2208,1302 $DEVICE_ID=1001
MM7 37 46 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2238 $Y=756  $PIN_XY=2268,672,2238,756,2208,672 $DEVICE_ID=1001
MM8 95 30 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=315  $PIN_XY=2268,378,2238,315,2208,378 $DEVICE_ID=1001
MM9 18 35 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1902 $Y=2243  $PIN_XY=1932,2226,1902,2243,1872,2226 $DEVICE_ID=1001
MM10 5 25 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=1197  $PIN_XY=1764,1302,1734,1197,1704,1302 $DEVICE_ID=1001
MM11 45 30 94 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=294  $PIN_XY=1764,378,1734,294,1704,378 $DEVICE_ID=1001
MM12 17 35 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1566 $Y=2244  $PIN_XY=1596,2226,1566,2244,1536,2226 $DEVICE_ID=1001
MM13 36 23 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1566 $Y=1680  $PIN_XY=1596,1596,1566,1680,1536,1596 $DEVICE_ID=1001
MM14 23 40 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=1218  $PIN_XY=1596,1302,1566,1218,1536,1302 $DEVICE_ID=1001
MM15 35 45 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1566 $Y=756  $PIN_XY=1596,672,1566,756,1536,672 $DEVICE_ID=1001
MM16 94 39 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=315  $PIN_XY=1596,378,1566,315,1536,378 $DEVICE_ID=1001
MM17 18 33 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1230 $Y=2243  $PIN_XY=1260,2226,1230,2243,1200,2226 $DEVICE_ID=1001
MM18 5 27 26 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=1197  $PIN_XY=1092,1302,1062,1197,1032,1302 $DEVICE_ID=1001
MM19 44 43 93 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=294  $PIN_XY=1092,378,1062,294,1032,378 $DEVICE_ID=1001
MM20 17 33 20 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=894 $Y=2244  $PIN_XY=924,2226,894,2244,864,2226 $DEVICE_ID=1001
MM21 34 26 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=894 $Y=1680  $PIN_XY=924,1596,894,1680,864,1596 $DEVICE_ID=1001
MM22 26 42 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=1218  $PIN_XY=924,1302,894,1218,864,1302 $DEVICE_ID=1001
MM23 33 44 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=894 $Y=756  $PIN_XY=924,672,894,756,864,672 $DEVICE_ID=1001
MM24 93 29 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=315  $PIN_XY=924,378,894,315,864,378 $DEVICE_ID=1001
MM25 18 31 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=558 $Y=2243  $PIN_XY=588,2226,558,2243,528,2226 $DEVICE_ID=1001
MM26 5 27 28 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=1197  $PIN_XY=420,1302,390,1197,360,1302 $DEVICE_ID=1001
MM27 41 29 92 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=294  $PIN_XY=420,378,390,294,360,378 $DEVICE_ID=1001
MM28 17 31 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=2267  $PIN_XY=252,2226,222,2267,192,2226 $DEVICE_ID=1001
MM29 32 28 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=1680  $PIN_XY=252,1596,222,1680,192,1596 $DEVICE_ID=1001
MM30 28 40 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=1218  $PIN_XY=252,1302,222,1218,192,1302 $DEVICE_ID=1001
MM31 31 41 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=756  $PIN_XY=252,672,222,756,192,672 $DEVICE_ID=1001
MM32 92 39 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=315  $PIN_XY=252,378,222,315,192,378 $DEVICE_ID=1001
MM33 6 24 38 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=1781  $PIN_XY=2436,1766,2406,1781,2376,1766 $DEVICE_ID=1003
MM34 24 25 88 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=1197  $PIN_XY=2436,1132,2406,1197,2376,1132 $DEVICE_ID=1003
MM35 4 46 37 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=857  $PIN_XY=2436,842,2406,857,2376,842 $DEVICE_ID=1003
MM36 38 24 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=1680  $PIN_XY=2268,1766,2238,1680,2208,1766 $DEVICE_ID=1003
MM37 88 42 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=1218  $PIN_XY=2268,1132,2238,1218,2208,1132 $DEVICE_ID=1003
MM38 37 46 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=756  $PIN_XY=2268,842,2238,756,2208,842 $DEVICE_ID=1003
MM39 6 23 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=1781  $PIN_XY=1764,1766,1734,1781,1704,1766 $DEVICE_ID=1003
MM40 23 25 89 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=1197  $PIN_XY=1764,1132,1734,1197,1704,1132 $DEVICE_ID=1003
MM41 4 45 35 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=857  $PIN_XY=1764,842,1734,857,1704,842 $DEVICE_ID=1003
MM42 36 23 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=1680  $PIN_XY=1596,1766,1566,1680,1536,1766 $DEVICE_ID=1003
MM43 89 40 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=1218  $PIN_XY=1596,1132,1566,1218,1536,1132 $DEVICE_ID=1003
MM44 35 45 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=756  $PIN_XY=1596,842,1566,756,1536,842 $DEVICE_ID=1003
MM45 6 26 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=1781  $PIN_XY=1092,1766,1062,1781,1032,1766 $DEVICE_ID=1003
MM46 26 27 90 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=1197  $PIN_XY=1092,1132,1062,1197,1032,1132 $DEVICE_ID=1003
MM47 4 44 33 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=857  $PIN_XY=1092,842,1062,857,1032,842 $DEVICE_ID=1003
MM48 34 26 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=1680  $PIN_XY=924,1766,894,1680,864,1766 $DEVICE_ID=1003
MM49 90 42 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=1218  $PIN_XY=924,1132,894,1218,864,1132 $DEVICE_ID=1003
MM50 33 44 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=756  $PIN_XY=924,842,894,756,864,842 $DEVICE_ID=1003
MM51 6 28 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=1781  $PIN_XY=420,1766,390,1781,360,1766 $DEVICE_ID=1003
MM52 28 27 91 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=1197  $PIN_XY=420,1132,390,1197,360,1132 $DEVICE_ID=1003
MM53 4 41 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=857  $PIN_XY=420,842,390,857,360,842 $DEVICE_ID=1003
MM54 32 28 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=1680  $PIN_XY=252,1766,222,1680,192,1766 $DEVICE_ID=1003
MM55 91 40 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=1218  $PIN_XY=252,1132,222,1218,192,1132 $DEVICE_ID=1003
MM56 31 41 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=756  $PIN_XY=252,842,222,756,192,842 $DEVICE_ID=1003
XX30BB92C5999 5 6 36 23 79 83 inv $T=1344 1386 0 0 $X=1344 $Y=1386
XX30BB92C51000 5 6 38 24 79 83 inv $T=2016 1386 0 0 $X=2016 $Y=1386
XX30BB92C51001 5 6 34 26 79 83 inv $T=672 1386 0 0 $X=672 $Y=1386
XX30BB92C51002 5 6 32 28 79 83 inv $T=0 1386 0 0 $X=0 $Y=1386
XX30BB92C51003 3 4 37 46 80 84 inv $T=2016 462 0 0 $X=2016 $Y=462
XX30BB92C51004 3 4 35 45 80 84 inv $T=1344 462 0 0 $X=1344 $Y=462
XX30BB92C51005 3 4 33 44 80 84 inv $T=672 462 0 0 $X=672 $Y=462
XX30BB92C51006 3 4 31 41 80 84 inv $T=0 462 0 0 $X=0 $Y=462
XX30BB92C51007 5 4 24 25 42 88 79 84 nor $T=1388 1514 1 0 $X=2016 $Y=922
XX30BB92C51008 5 4 23 25 40 89 79 84 nor $T=716 1514 1 0 $X=1343 $Y=922
XX30BB92C51009 5 4 26 27 42 90 79 84 nor $T=44 1514 1 0 $X=672 $Y=922
XX30BB92C51010 5 4 28 27 40 91 79 84 nor $T=-628 1514 1 0 $X=0 $Y=922
XX30BB92C51011 3 2 41 39 29 92 80 85 nand $T=-418 816 1 0 $X=0 $Y=-2
XX30BB92C51012 3 2 44 29 43 93 80 85 nand $T=254 816 1 0 $X=671 $Y=-2
XX30BB92C51013 3 2 45 39 30 94 80 85 nand $T=926 816 1 0 $X=1344 $Y=-2
XX30BB92C51014 3 2 46 30 43 95 80 85 nand $T=1598 816 1 0 $X=2016 $Y=-2
.ends 2to4_decoder_static
.subckt between_blocks 2 3 4 5 6 7 8 9 10 12 13
+	15 16 17 18 19 20 25 26 27 28 29
+	30 31 32 33 34 35 36 37 38 39 40
+	41 42 43 44 53
MM1 9 22 28 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1390 $Y=1777  $PIN_XY=1420,1882,1390,1777,1360,1882 $DEVICE_ID=1001
MM2 7 21 34 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1390 $Y=853  $PIN_XY=1420,958,1390,853,1360,958 $DEVICE_ID=1001
MM3 5 14 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1390 $Y=-71  $PIN_XY=1420,34,1390,-71,1360,34 $DEVICE_ID=1001
MM4 2 13 30 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1390 $Y=-974  $PIN_XY=1420,-890,1390,-974,1360,-890 $DEVICE_ID=1001
MM5 35 12 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1222 $Y=2260  $PIN_XY=1252,2176,1222,2260,1192,2176 $DEVICE_ID=1001
MM6 29 11 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1222 $Y=1357  $PIN_XY=1252,1252,1222,1357,1192,1252 $DEVICE_ID=1001
MM7 45 24 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1222 $Y=433  $PIN_XY=1252,328,1222,433,1192,328 $DEVICE_ID=1001
MM8 31 23 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1222 $Y=-491  $PIN_XY=1252,-596,1222,-491,1192,-596 $DEVICE_ID=1001
MM9 9 15 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=1798  $PIN_XY=916,1882,886,1798,856,1882 $DEVICE_ID=1001
MM10 7 15 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=874  $PIN_XY=916,958,886,874,856,958 $DEVICE_ID=1001
MM11 5 32 51 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=-50  $PIN_XY=916,34,886,-50,856,34 $DEVICE_ID=1001
MM12 2 16 49 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=-974  $PIN_XY=916,-890,886,-974,856,-890 $DEVICE_ID=1001
MM13 9 19 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=2239  $PIN_XY=748,2176,718,2239,688,2176 $DEVICE_ID=1001
MM14 22 20 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=1798  $PIN_XY=748,1882,718,1798,688,1882 $DEVICE_ID=1001
MM15 7 18 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=1336  $PIN_XY=748,1252,718,1336,688,1252 $DEVICE_ID=1001
MM16 21 17 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=874  $PIN_XY=748,958,718,874,688,958 $DEVICE_ID=1001
MM17 24 27 52 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=412  $PIN_XY=748,328,718,412,688,328 $DEVICE_ID=1001
MM18 51 16 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=-50  $PIN_XY=748,34,718,-50,688,34 $DEVICE_ID=1001
MM19 23 26 50 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=-512  $PIN_XY=748,-596,718,-512,688,-596 $DEVICE_ID=1001
MM20 49 25 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=-953  $PIN_XY=748,-890,718,-953,688,-890 $DEVICE_ID=1001
MM21 12 15 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=2260  $PIN_XY=580,2176,550,2260,520,2176 $DEVICE_ID=1001
MM22 11 15 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=1336  $PIN_XY=580,1252,550,1336,520,1252 $DEVICE_ID=1001
MM23 52 16 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=412  $PIN_XY=580,328,550,412,520,328 $DEVICE_ID=1001
MM24 50 16 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=-512  $PIN_XY=580,-596,550,-512,520,-596 $DEVICE_ID=1001
MM25 8 22 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=1777  $PIN_XY=1420,1712,1390,1777,1360,1712 $DEVICE_ID=1003
MM26 8 11 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=1437  $PIN_XY=1420,1422,1390,1437,1360,1422 $DEVICE_ID=1003
MM27 6 21 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=853  $PIN_XY=1420,788,1390,853,1360,788 $DEVICE_ID=1003
MM28 6 24 45 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=513  $PIN_XY=1420,498,1390,513,1360,498 $DEVICE_ID=1003
MM29 4 14 33 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=-71  $PIN_XY=1420,-136,1390,-71,1360,-136 $DEVICE_ID=1003
MM30 4 23 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=-411  $PIN_XY=1420,-426,1390,-411,1360,-426 $DEVICE_ID=1003
MM31 28 22 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=1697  $PIN_XY=1252,1712,1222,1697,1192,1712 $DEVICE_ID=1003
MM32 29 11 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=1357  $PIN_XY=1252,1422,1222,1357,1192,1422 $DEVICE_ID=1003
MM33 34 21 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=773  $PIN_XY=1252,788,1222,773,1192,788 $DEVICE_ID=1003
MM34 45 24 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=433  $PIN_XY=1252,498,1222,433,1192,498 $DEVICE_ID=1003
MM35 33 14 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=-151  $PIN_XY=1252,-136,1222,-151,1192,-136 $DEVICE_ID=1003
MM36 31 23 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=-491  $PIN_XY=1252,-426,1222,-491,1192,-426 $DEVICE_ID=1003
MM37 8 15 48 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=1798  $PIN_XY=916,1712,886,1798,856,1712 $DEVICE_ID=1003
MM38 6 15 46 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=874  $PIN_XY=916,788,886,874,856,788 $DEVICE_ID=1003
MM39 4 32 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=-50  $PIN_XY=916,-136,886,-50,856,-136 $DEVICE_ID=1003
MM40 48 20 22 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=1798  $PIN_XY=748,1712,718,1798,688,1712 $DEVICE_ID=1003
MM41 11 18 47 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=1336  $PIN_XY=748,1422,718,1336,688,1422 $DEVICE_ID=1003
MM42 46 17 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=874  $PIN_XY=748,788,718,874,688,788 $DEVICE_ID=1003
MM43 6 27 24 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=412  $PIN_XY=748,498,718,412,688,498 $DEVICE_ID=1003
MM44 14 16 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=-50  $PIN_XY=748,-136,718,-50,688,-136 $DEVICE_ID=1003
MM45 4 26 23 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=-512  $PIN_XY=748,-426,718,-512,688,-426 $DEVICE_ID=1003
MM46 47 15 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=1336  $PIN_XY=580,1422,550,1336,520,1422 $DEVICE_ID=1003
MM47 24 16 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=412  $PIN_XY=580,498,550,412,520,498 $DEVICE_ID=1003
MM48 23 16 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=-512  $PIN_XY=580,-426,550,-512,520,-426 $DEVICE_ID=1003
XX30BB92C51015 2 3 30 13 36 40 inv $T=1612 -680 0 180 $X=1000 $Y=-1270
XX30BB92C51016 2 4 31 23 36 41 inv $T=1000 -806 0 0 $X=1000 $Y=-806
XX30BB92C51017 5 4 33 14 37 41 inv $T=1612 244 0 180 $X=1000 $Y=-346
XX30BB92C51018 5 6 45 24 37 42 inv $T=1000 118 0 0 $X=1000 $Y=118
XX30BB92C51019 7 6 34 21 38 42 inv $T=1612 1168 0 180 $X=1000 $Y=578
XX30BB92C51020 7 8 29 11 38 43 inv $T=1000 1042 0 0 $X=1000 $Y=1042
XX30BB92C51021 9 8 28 22 39 43 inv $T=1612 2092 0 180 $X=1000 $Y=1502
XX30BB92C51022 9 10 35 12 39 44 inv $T=1000 1966 0 0 $X=1000 $Y=1966
XX30BB92C51023 7 6 21 17 15 46 38 42 nor $T=1736 1170 0 180 $X=328 $Y=578
XX30BB92C51024 7 8 11 18 15 47 38 43 nor $T=-300 1040 0 0 $X=328 $Y=1042
XX30BB92C51025 9 8 22 20 15 48 39 43 nor $T=1736 2094 0 180 $X=328 $Y=1501
XX30BB92C51026 9 10 12 19 15 53 39 44 nor $T=-300 1964 0 0 $X=328 $Y=1966
XX30BB92C51027 2 3 13 16 25 49 36 40 nand $T=1526 -452 0 180 $X=328 $Y=-1270
XX30BB92C51028 2 4 23 16 26 50 36 41 nand $T=-90 -1034 0 0 $X=327 $Y=-806
XX30BB92C51029 5 4 14 32 16 51 37 41 nand $T=1526 472 0 180 $X=328 $Y=-346
XX30BB92C51030 5 6 24 16 27 52 37 42 nand $T=-90 -110 0 0 $X=327 $Y=118
.ends between_blocks
.subckt read_circuit 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16
XX30BB92C51040 2 3 5 4 14 15 invx4 $T=-24 4 0 0 $X=0 $Y=4
XX30BB92C51041 2 3 8 7 14 15 inv $T=1512 4 0 0 $X=1512 $Y=4
XX30BB92C51042 2 3 7 5 6 16 14 15 nand $T=422 -224 0 0 $X=840 $Y=4
.ends read_circuit
.subckt buffer_highdrive 2 3 4 5 6 7 8 9
XX30BB92C51043 3 2 5 6 8 9 invx4 $T=-22 -2 0 0 $X=2 $Y=-2
XX30BB92C51044 3 2 4 5 8 9 invx4 $T=818 -2 0 0 $X=842 $Y=-2
.ends buffer_highdrive
.subckt buffer 2 3 4 5 6 7 8
XX30BB92C51045 2 3 5 4 7 8 inv $T=584 2 0 0 $X=584 $Y=2
XX30BB92C51046 2 3 4 6 7 8 inv $T=80 2 0 0 $X=80 $Y=2
.ends buffer
.subckt Demux 2 3 4 5 6 7 8 9 10 11 12
+	13 14
MM1 11 9 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1398 $Y=735  $PIN_XY=1428,672,1398,735,1368,672 $DEVICE_ID=1001
MM2 10 8 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1398 $Y=315  $PIN_XY=1428,378,1398,315,1368,378 $DEVICE_ID=1001
MM3 9 6 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=894 $Y=735  $PIN_XY=924,672,894,735,864,672 $DEVICE_ID=1001
MM4 8 5 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=894 $Y=315  $PIN_XY=924,378,894,315,864,378 $DEVICE_ID=1001
MM5 15 7 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=726 $Y=735  $PIN_XY=756,672,726,735,696,672 $DEVICE_ID=1001
MM6 16 7 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=726 $Y=315  $PIN_XY=756,378,726,315,696,378 $DEVICE_ID=1001
MM7 6 5 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=756  $PIN_XY=252,672,222,756,192,672 $DEVICE_ID=1001
XX30BB92C51047 2 3 _GENERATED_17 2 12 13 sram_filler $T=616 588 0 180 $X=167 $Y=-2
XX30BB92C51048 2 3 3 _GENERATED_18 12 13 sram_filler $T=448 588 0 180 $X=0 $Y=-2
XX30BB92C51049 2 4 6 5 12 14 inv $T=0 462 0 0 $X=0 $Y=462
XX30BB92C51050 2 4 11 9 12 14 inv $T=1176 462 0 0 $X=1176 $Y=462
XX30BB92C51051 2 3 10 8 12 13 inv $T=1176 588 1 0 $X=1176 $Y=-2
XX30BB92C51052 2 4 9 7 6 15 12 14 nand $T=86 234 0 0 $X=504 $Y=462
XX30BB92C51053 2 3 8 7 5 16 12 13 nand $T=86 816 1 0 $X=504 $Y=-2
.ends Demux

* Hierarchy Level 1
.subckt static_row_decoder_3by8 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16 17 18 26 27 28 31 32
+	34 51 52 53 54 55 56 57 58 59 60
+	61 62 63 64 65 66 67 68 69 70 71
+	72 73 74 75 88 112
*.floating_nets 107 108 109 110 111
MM1 16 90 57 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=884  $PIN_XY=3760,800,3730,884,3700,800 $DEVICE_ID=1001
MM2 11 91 58 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-40  $PIN_XY=3760,-124,3730,-40,3700,-124 $DEVICE_ID=1001
MM3 10 87 54 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-964  $PIN_XY=3760,-1048,3730,-964,3700,-1048 $DEVICE_ID=1001
MM4 13 86 53 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-1888  $PIN_XY=3760,-1972,3730,-1888,3700,-1972 $DEVICE_ID=1001
MM5 5 84 51 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-2812  $PIN_XY=3760,-2896,3730,-2812,3700,-2896 $DEVICE_ID=1001
MM6 8 89 56 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-3736  $PIN_XY=3760,-3820,3730,-3736,3700,-3820 $DEVICE_ID=1001
MM7 3 85 52 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-4660  $PIN_XY=3760,-4744,3730,-4660,3700,-4744 $DEVICE_ID=1001
MM8 57 90 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=884  $PIN_XY=3592,800,3562,884,3532,800 $DEVICE_ID=1001
MM9 58 91 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-40  $PIN_XY=3592,-124,3562,-40,3532,-124 $DEVICE_ID=1001
MM10 54 87 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-964  $PIN_XY=3592,-1048,3562,-964,3532,-1048 $DEVICE_ID=1001
MM11 53 86 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-1888  $PIN_XY=3592,-1972,3562,-1888,3532,-1972 $DEVICE_ID=1001
MM12 51 84 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-2812  $PIN_XY=3592,-2896,3562,-2812,3532,-2896 $DEVICE_ID=1001
MM13 56 89 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-3736  $PIN_XY=3592,-3820,3562,-3736,3532,-3820 $DEVICE_ID=1001
MM14 52 85 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-4660  $PIN_XY=3592,-4744,3562,-4660,3532,-4744 $DEVICE_ID=1001
MM15 15 50 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=1346  $PIN_XY=2920,1430,2890,1346,2860,1430 $DEVICE_ID=1001
MM16 16 25 90 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=884  $PIN_XY=2920,800,2890,884,2860,800 $DEVICE_ID=1001
MM17 16 49 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=422  $PIN_XY=2920,506,2890,422,2860,506 $DEVICE_ID=1001
MM18 11 24 91 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-40  $PIN_XY=2920,-124,2890,-40,2860,-124 $DEVICE_ID=1001
MM19 11 48 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-502  $PIN_XY=2920,-418,2890,-502,2860,-418 $DEVICE_ID=1001
MM20 10 23 87 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-964  $PIN_XY=2920,-1048,2890,-964,2860,-1048 $DEVICE_ID=1001
MM21 10 47 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-1426  $PIN_XY=2920,-1342,2890,-1426,2860,-1342 $DEVICE_ID=1001
MM22 13 22 86 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-1888  $PIN_XY=2920,-1972,2890,-1888,2860,-1972 $DEVICE_ID=1001
MM23 13 43 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-2350  $PIN_XY=2920,-2266,2890,-2350,2860,-2266 $DEVICE_ID=1001
MM24 5 21 84 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-2812  $PIN_XY=2920,-2896,2890,-2812,2860,-2896 $DEVICE_ID=1001
MM25 5 42 20 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-3274  $PIN_XY=2920,-3190,2890,-3274,2860,-3190 $DEVICE_ID=1001
MM26 8 20 89 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-3736  $PIN_XY=2920,-3820,2890,-3736,2860,-3820 $DEVICE_ID=1001
MM27 8 41 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-4198  $PIN_XY=2920,-4114,2890,-4198,2860,-4114 $DEVICE_ID=1001
MM28 3 19 85 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-4660  $PIN_XY=2920,-4744,2890,-4660,2860,-4744 $DEVICE_ID=1001
MM29 25 46 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=1346  $PIN_XY=2752,1430,2722,1346,2692,1430 $DEVICE_ID=1001
MM30 90 25 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=884  $PIN_XY=2752,800,2722,884,2692,800 $DEVICE_ID=1001
MM31 24 45 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=422  $PIN_XY=2752,506,2722,422,2692,506 $DEVICE_ID=1001
MM32 91 24 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-40  $PIN_XY=2752,-124,2722,-40,2692,-124 $DEVICE_ID=1001
MM33 23 44 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-502  $PIN_XY=2752,-418,2722,-502,2692,-418 $DEVICE_ID=1001
MM34 87 23 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-964  $PIN_XY=2752,-1048,2722,-964,2692,-1048 $DEVICE_ID=1001
MM35 22 40 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-1426  $PIN_XY=2752,-1342,2722,-1426,2692,-1342 $DEVICE_ID=1001
MM36 86 22 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-1888  $PIN_XY=2752,-1972,2722,-1888,2692,-1972 $DEVICE_ID=1001
MM37 21 39 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-2350  $PIN_XY=2752,-2266,2722,-2350,2692,-2266 $DEVICE_ID=1001
MM38 84 21 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-2812  $PIN_XY=2752,-2896,2722,-2812,2692,-2896 $DEVICE_ID=1001
MM39 20 38 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-3274  $PIN_XY=2752,-3190,2722,-3274,2692,-3190 $DEVICE_ID=1001
MM40 89 20 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-3736  $PIN_XY=2752,-3820,2722,-3736,2692,-3820 $DEVICE_ID=1001
MM41 19 37 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-4198  $PIN_XY=2752,-4114,2722,-4198,2692,-4114 $DEVICE_ID=1001
MM42 85 19 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-4660  $PIN_XY=2752,-4744,2722,-4660,2692,-4744 $DEVICE_ID=1001
MM43 50 36 105 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=1346  $PIN_XY=2248,1430,2218,1346,2188,1430 $DEVICE_ID=1001
MM44 46 28 106 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=884  $PIN_XY=2248,800,2218,884,2188,800 $DEVICE_ID=1001
MM45 49 36 104 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=422  $PIN_XY=2248,506,2218,422,2188,506 $DEVICE_ID=1001
MM46 45 28 99 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-40  $PIN_XY=2248,-124,2218,-40,2188,-124 $DEVICE_ID=1001
MM47 48 27 102 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-502  $PIN_XY=2248,-418,2218,-502,2188,-418 $DEVICE_ID=1001
MM48 44 28 103 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-964  $PIN_XY=2248,-1048,2218,-964,2188,-1048 $DEVICE_ID=1001
MM49 47 27 101 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-1426  $PIN_XY=2248,-1342,2218,-1426,2188,-1342 $DEVICE_ID=1001
MM50 40 28 100 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-1888  $PIN_XY=2248,-1972,2218,-1888,2188,-1972 $DEVICE_ID=1001
MM51 43 36 93 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-2350  $PIN_XY=2248,-2266,2218,-2350,2188,-2266 $DEVICE_ID=1001
MM52 39 28 92 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-2812  $PIN_XY=2248,-2896,2218,-2812,2188,-2896 $DEVICE_ID=1001
MM53 42 36 94 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-3274  $PIN_XY=2248,-3190,2218,-3274,2188,-3190 $DEVICE_ID=1001
MM54 38 28 95 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-3736  $PIN_XY=2248,-3820,2218,-3736,2188,-3820 $DEVICE_ID=1001
MM55 41 27 97 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-4198  $PIN_XY=2248,-4114,2218,-4198,2188,-4114 $DEVICE_ID=1001
MM56 37 28 96 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-4660  $PIN_XY=2248,-4744,2218,-4660,2188,-4744 $DEVICE_ID=1001
MM57 105 29 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=1346  $PIN_XY=2080,1430,2050,1346,2020,1430 $DEVICE_ID=1001
MM58 106 35 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=884  $PIN_XY=2080,800,2050,884,2020,800 $DEVICE_ID=1001
MM59 104 26 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=422  $PIN_XY=2080,506,2050,422,2020,506 $DEVICE_ID=1001
MM60 99 35 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-40  $PIN_XY=2080,-124,2050,-40,2020,-124 $DEVICE_ID=1001
MM61 102 29 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-502  $PIN_XY=2080,-418,2050,-502,2020,-418 $DEVICE_ID=1001
MM62 103 35 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-964  $PIN_XY=2080,-1048,2050,-964,2020,-1048 $DEVICE_ID=1001
MM63 101 26 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-1426  $PIN_XY=2080,-1342,2050,-1426,2020,-1342 $DEVICE_ID=1001
MM64 100 35 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-1888  $PIN_XY=2080,-1972,2050,-1888,2020,-1972 $DEVICE_ID=1001
MM65 93 29 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-2350  $PIN_XY=2080,-2266,2050,-2350,2020,-2266 $DEVICE_ID=1001
MM66 92 31 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-2812  $PIN_XY=2080,-2896,2050,-2812,2020,-2896 $DEVICE_ID=1001
MM67 94 31 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-3274  $PIN_XY=2080,-3190,2050,-3274,2020,-3190 $DEVICE_ID=1001
MM68 95 26 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-3736  $PIN_XY=2080,-3820,2050,-3736,2020,-3820 $DEVICE_ID=1001
MM69 97 29 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-4198  $PIN_XY=2080,-4114,2050,-4198,2020,-4114 $DEVICE_ID=1001
MM70 96 31 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-4660  $PIN_XY=2080,-4744,2050,-4660,2020,-4744 $DEVICE_ID=1001
MM71 29 26 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1546 $Y=1346  $PIN_XY=1576,1430,1546,1346,1516,1430 $DEVICE_ID=1001
MM72 36 27 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1546 $Y=884  $PIN_XY=1576,800,1546,884,1516,800 $DEVICE_ID=1001
MM73 35 31 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1546 $Y=443  $PIN_XY=1576,506,1546,443,1516,506 $DEVICE_ID=1001
MM74 3 34 30 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1042 $Y=-4681  $PIN_XY=1072,-4744,1042,-4681,1012,-4744 $DEVICE_ID=1001
MM75 30 34 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=874 $Y=-4681  $PIN_XY=904,-4744,874,-4681,844,-4744 $DEVICE_ID=1001
MM76 3 33 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-5122  $PIN_XY=2920,-5038,2890,-5122,2860,-5038 $DEVICE_ID=1001
MM77 18 32 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-5122  $PIN_XY=2752,-5038,2722,-5122,2692,-5038 $DEVICE_ID=1001
MM78 33 27 98 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-5122  $PIN_XY=2248,-5038,2218,-5122,2188,-5038 $DEVICE_ID=1001
MM79 98 31 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-5122  $PIN_XY=2080,-5038,2050,-5122,2020,-5038 $DEVICE_ID=1001
MM80 3 30 28 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1042 $Y=-5101  $PIN_XY=1072,-5038,1042,-5101,1012,-5038 $DEVICE_ID=1001
MM81 28 30 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=874 $Y=-5101  $PIN_XY=904,-5038,874,-5101,844,-5038 $DEVICE_ID=1001
MM82 14 90 57 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=964  $PIN_XY=4096,970,4066,964,4036,970 $DEVICE_ID=1003
MM83 17 91 58 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=40  $PIN_XY=4096,46,4066,40,4036,46 $DEVICE_ID=1003
MM84 9 87 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-884  $PIN_XY=4096,-878,4066,-884,4036,-878 $DEVICE_ID=1003
MM85 12 86 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-1808  $PIN_XY=4096,-1802,4066,-1808,4036,-1802 $DEVICE_ID=1003
MM86 6 84 51 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-2732  $PIN_XY=4096,-2726,4066,-2732,4036,-2726 $DEVICE_ID=1003
MM87 7 89 56 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-3656  $PIN_XY=4096,-3650,4066,-3656,4036,-3650 $DEVICE_ID=1003
MM88 2 85 52 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-4580  $PIN_XY=4096,-4574,4066,-4580,4036,-4574 $DEVICE_ID=1003
MM89 57 90 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=964  $PIN_XY=3928,970,3898,964,3868,970 $DEVICE_ID=1003
MM90 58 91 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=40  $PIN_XY=3928,46,3898,40,3868,46 $DEVICE_ID=1003
MM91 54 87 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-884  $PIN_XY=3928,-878,3898,-884,3868,-878 $DEVICE_ID=1003
MM92 53 86 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-1808  $PIN_XY=3928,-1802,3898,-1808,3868,-1802 $DEVICE_ID=1003
MM93 51 84 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-2732  $PIN_XY=3928,-2726,3898,-2732,3868,-2726 $DEVICE_ID=1003
MM94 56 89 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-3656  $PIN_XY=3928,-3650,3898,-3656,3868,-3650 $DEVICE_ID=1003
MM95 52 85 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-4580  $PIN_XY=3928,-4574,3898,-4580,3868,-4574 $DEVICE_ID=1003
MM96 14 90 57 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=884  $PIN_XY=3760,970,3730,884,3700,970 $DEVICE_ID=1003
MM97 17 91 58 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-40  $PIN_XY=3760,46,3730,-40,3700,46 $DEVICE_ID=1003
MM98 9 87 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-964  $PIN_XY=3760,-878,3730,-964,3700,-878 $DEVICE_ID=1003
MM99 12 86 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-1888  $PIN_XY=3760,-1802,3730,-1888,3700,-1802 $DEVICE_ID=1003
MM100 6 84 51 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-2812  $PIN_XY=3760,-2726,3730,-2812,3700,-2726 $DEVICE_ID=1003
MM101 7 89 56 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-3736  $PIN_XY=3760,-3650,3730,-3736,3700,-3650 $DEVICE_ID=1003
MM102 57 90 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=884  $PIN_XY=3592,970,3562,884,3532,970 $DEVICE_ID=1003
MM103 58 91 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-40  $PIN_XY=3592,46,3562,-40,3532,46 $DEVICE_ID=1003
MM104 54 87 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-964  $PIN_XY=3592,-878,3562,-964,3532,-878 $DEVICE_ID=1003
MM105 53 86 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-1888  $PIN_XY=3592,-1802,3562,-1888,3532,-1802 $DEVICE_ID=1003
MM106 51 84 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-2812  $PIN_XY=3592,-2726,3562,-2812,3532,-2726 $DEVICE_ID=1003
MM107 56 89 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-3736  $PIN_XY=3592,-3650,3562,-3736,3532,-3650 $DEVICE_ID=1003
MM108 14 25 90 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=964  $PIN_XY=3256,970,3226,964,3196,970 $DEVICE_ID=1003
MM109 17 24 91 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=40  $PIN_XY=3256,46,3226,40,3196,46 $DEVICE_ID=1003
MM110 9 23 87 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-884  $PIN_XY=3256,-878,3226,-884,3196,-878 $DEVICE_ID=1003
MM111 12 22 86 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-1808  $PIN_XY=3256,-1802,3226,-1808,3196,-1802 $DEVICE_ID=1003
MM112 6 21 84 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-2732  $PIN_XY=3256,-2726,3226,-2732,3196,-2726 $DEVICE_ID=1003
MM113 7 20 89 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-3656  $PIN_XY=3256,-3650,3226,-3656,3196,-3650 $DEVICE_ID=1003
MM114 2 19 85 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-4580  $PIN_XY=3256,-4574,3226,-4580,3196,-4574 $DEVICE_ID=1003
MM115 90 25 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=964  $PIN_XY=3088,970,3058,964,3028,970 $DEVICE_ID=1003
MM116 91 24 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=40  $PIN_XY=3088,46,3058,40,3028,46 $DEVICE_ID=1003
MM117 87 23 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-884  $PIN_XY=3088,-878,3058,-884,3028,-878 $DEVICE_ID=1003
MM118 86 22 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-1808  $PIN_XY=3088,-1802,3058,-1808,3028,-1802 $DEVICE_ID=1003
MM119 84 21 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-2732  $PIN_XY=3088,-2726,3058,-2732,3028,-2726 $DEVICE_ID=1003
MM120 89 20 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-3656  $PIN_XY=3088,-3650,3058,-3656,3028,-3650 $DEVICE_ID=1003
MM121 85 19 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-4580  $PIN_XY=3088,-4574,3058,-4580,3028,-4574 $DEVICE_ID=1003
MM122 25 50 82 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=1346  $PIN_XY=2920,1260,2890,1346,2860,1260 $DEVICE_ID=1003
MM123 14 25 90 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=884  $PIN_XY=2920,970,2890,884,2860,970 $DEVICE_ID=1003
MM124 24 49 83 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=422  $PIN_XY=2920,336,2890,422,2860,336 $DEVICE_ID=1003
MM125 17 24 91 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-40  $PIN_XY=2920,46,2890,-40,2860,46 $DEVICE_ID=1003
MM126 23 48 81 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-502  $PIN_XY=2920,-588,2890,-502,2860,-588 $DEVICE_ID=1003
MM127 9 23 87 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-964  $PIN_XY=2920,-878,2890,-964,2860,-878 $DEVICE_ID=1003
MM128 22 47 80 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-1426  $PIN_XY=2920,-1512,2890,-1426,2860,-1512 $DEVICE_ID=1003
MM129 12 22 86 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-1888  $PIN_XY=2920,-1802,2890,-1888,2860,-1802 $DEVICE_ID=1003
MM130 21 43 77 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-2350  $PIN_XY=2920,-2436,2890,-2350,2860,-2436 $DEVICE_ID=1003
MM131 6 21 84 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-2812  $PIN_XY=2920,-2726,2890,-2812,2860,-2726 $DEVICE_ID=1003
MM132 20 42 78 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-3274  $PIN_XY=2920,-3360,2890,-3274,2860,-3360 $DEVICE_ID=1003
MM133 7 20 89 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-3736  $PIN_XY=2920,-3650,2890,-3736,2860,-3650 $DEVICE_ID=1003
MM134 19 41 76 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-4198  $PIN_XY=2920,-4284,2890,-4198,2860,-4284 $DEVICE_ID=1003
MM135 82 46 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=1346  $PIN_XY=2752,1260,2722,1346,2692,1260 $DEVICE_ID=1003
MM136 90 25 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=884  $PIN_XY=2752,970,2722,884,2692,970 $DEVICE_ID=1003
MM137 83 45 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=422  $PIN_XY=2752,336,2722,422,2692,336 $DEVICE_ID=1003
MM138 91 24 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-40  $PIN_XY=2752,46,2722,-40,2692,46 $DEVICE_ID=1003
MM139 81 44 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-502  $PIN_XY=2752,-588,2722,-502,2692,-588 $DEVICE_ID=1003
MM140 87 23 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-964  $PIN_XY=2752,-878,2722,-964,2692,-878 $DEVICE_ID=1003
MM141 80 40 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-1426  $PIN_XY=2752,-1512,2722,-1426,2692,-1512 $DEVICE_ID=1003
MM142 86 22 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-1888  $PIN_XY=2752,-1802,2722,-1888,2692,-1802 $DEVICE_ID=1003
MM143 77 39 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-2350  $PIN_XY=2752,-2436,2722,-2350,2692,-2436 $DEVICE_ID=1003
MM144 84 21 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-2812  $PIN_XY=2752,-2726,2722,-2812,2692,-2726 $DEVICE_ID=1003
MM145 78 38 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-3274  $PIN_XY=2752,-3360,2722,-3274,2692,-3360 $DEVICE_ID=1003
MM146 89 20 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-3736  $PIN_XY=2752,-3650,2722,-3736,2692,-3650 $DEVICE_ID=1003
MM147 76 37 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-4198  $PIN_XY=2752,-4284,2722,-4198,2692,-4284 $DEVICE_ID=1003
MM148 14 36 50 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=1346  $PIN_XY=2248,1260,2218,1346,2188,1260 $DEVICE_ID=1003
MM149 14 28 46 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=884  $PIN_XY=2248,970,2218,884,2188,970 $DEVICE_ID=1003
MM150 17 36 49 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=422  $PIN_XY=2248,336,2218,422,2188,336 $DEVICE_ID=1003
MM151 17 28 45 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-40  $PIN_XY=2248,46,2218,-40,2188,46 $DEVICE_ID=1003
MM152 9 27 48 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-502  $PIN_XY=2248,-588,2218,-502,2188,-588 $DEVICE_ID=1003
MM153 9 28 44 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-964  $PIN_XY=2248,-878,2218,-964,2188,-878 $DEVICE_ID=1003
MM154 12 27 47 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-1426  $PIN_XY=2248,-1512,2218,-1426,2188,-1512 $DEVICE_ID=1003
MM155 12 28 40 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-1888  $PIN_XY=2248,-1802,2218,-1888,2188,-1802 $DEVICE_ID=1003
MM156 6 36 43 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-2350  $PIN_XY=2248,-2436,2218,-2350,2188,-2436 $DEVICE_ID=1003
MM157 6 28 39 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-2812  $PIN_XY=2248,-2726,2218,-2812,2188,-2726 $DEVICE_ID=1003
MM158 7 36 42 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-3274  $PIN_XY=2248,-3360,2218,-3274,2188,-3360 $DEVICE_ID=1003
MM159 7 28 38 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-3736  $PIN_XY=2248,-3650,2218,-3736,2188,-3650 $DEVICE_ID=1003
MM160 2 27 41 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-4198  $PIN_XY=2248,-4284,2218,-4198,2188,-4284 $DEVICE_ID=1003
MM161 50 29 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=1346  $PIN_XY=2080,1260,2050,1346,2020,1260 $DEVICE_ID=1003
MM162 46 35 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=884  $PIN_XY=2080,970,2050,884,2020,970 $DEVICE_ID=1003
MM163 49 26 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=422  $PIN_XY=2080,336,2050,422,2020,336 $DEVICE_ID=1003
MM164 45 35 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-40  $PIN_XY=2080,46,2050,-40,2020,46 $DEVICE_ID=1003
MM165 48 29 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-502  $PIN_XY=2080,-588,2050,-502,2020,-588 $DEVICE_ID=1003
MM166 44 35 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-964  $PIN_XY=2080,-878,2050,-964,2020,-878 $DEVICE_ID=1003
MM167 47 26 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-1426  $PIN_XY=2080,-1512,2050,-1426,2020,-1512 $DEVICE_ID=1003
MM168 40 35 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-1888  $PIN_XY=2080,-1802,2050,-1888,2020,-1802 $DEVICE_ID=1003
MM169 43 29 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-2350  $PIN_XY=2080,-2436,2050,-2350,2020,-2436 $DEVICE_ID=1003
MM170 39 31 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-2812  $PIN_XY=2080,-2726,2050,-2812,2020,-2726 $DEVICE_ID=1003
MM171 42 31 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-3274  $PIN_XY=2080,-3360,2050,-3274,2020,-3360 $DEVICE_ID=1003
MM172 38 26 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-3736  $PIN_XY=2080,-3650,2050,-3736,2020,-3650 $DEVICE_ID=1003
MM173 41 29 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-4198  $PIN_XY=2080,-4284,2050,-4198,2020,-4284 $DEVICE_ID=1003
MM174 14 26 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1714 $Y=1245  $PIN_XY=1744,1260,1714,1245,1684,1260 $DEVICE_ID=1003
MM175 14 27 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1714 $Y=985  $PIN_XY=1744,970,1714,985,1684,970 $DEVICE_ID=1003
MM176 17 31 35 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1714 $Y=342  $PIN_XY=1744,336,1714,342,1684,336 $DEVICE_ID=1003
MM177 29 26 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1546 $Y=1346  $PIN_XY=1576,1260,1546,1346,1516,1260 $DEVICE_ID=1003
MM178 36 27 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1546 $Y=884  $PIN_XY=1576,970,1546,884,1516,970 $DEVICE_ID=1003
MM179 35 31 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1546 $Y=443  $PIN_XY=1576,336,1546,443,1516,336 $DEVICE_ID=1003
MM180 2 34 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1378 $Y=-4580  $PIN_XY=1408,-4574,1378,-4580,1348,-4574 $DEVICE_ID=1003
MM181 30 34 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1210 $Y=-4580  $PIN_XY=1240,-4574,1210,-4580,1180,-4574 $DEVICE_ID=1003
MM182 2 88 55 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-5504  $PIN_XY=4096,-5498,4066,-5504,4036,-5498 $DEVICE_ID=1003
MM183 55 88 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-5504  $PIN_XY=3928,-5498,3898,-5504,3868,-5498 $DEVICE_ID=1003
MM184 2 85 52 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-4660  $PIN_XY=3760,-4574,3730,-4660,3700,-4574 $DEVICE_ID=1003
MM185 2 88 55 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-5584  $PIN_XY=3760,-5498,3730,-5584,3700,-5498 $DEVICE_ID=1003
MM186 52 85 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-4660  $PIN_XY=3592,-4574,3562,-4660,3532,-4574 $DEVICE_ID=1003
MM187 55 88 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-5584  $PIN_XY=3592,-5498,3562,-5584,3532,-5498 $DEVICE_ID=1003
MM188 2 18 88 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-5504  $PIN_XY=3256,-5498,3226,-5504,3196,-5498 $DEVICE_ID=1003
MM189 88 18 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-5504  $PIN_XY=3088,-5498,3058,-5504,3028,-5498 $DEVICE_ID=1003
MM190 2 19 85 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-4660  $PIN_XY=2920,-4574,2890,-4660,2860,-4574 $DEVICE_ID=1003
MM191 18 33 79 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-5122  $PIN_XY=2920,-5208,2890,-5122,2860,-5208 $DEVICE_ID=1003
MM192 2 18 88 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-5563  $PIN_XY=2920,-5498,2890,-5563,2860,-5498 $DEVICE_ID=1003
MM193 85 19 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-4660  $PIN_XY=2752,-4574,2722,-4660,2692,-4574 $DEVICE_ID=1003
MM194 79 32 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-5122  $PIN_XY=2752,-5208,2722,-5122,2692,-5208 $DEVICE_ID=1003
MM195 88 18 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-5563  $PIN_XY=2752,-5498,2722,-5563,2692,-5498 $DEVICE_ID=1003
MM196 2 28 37 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-4660  $PIN_XY=2248,-4574,2218,-4660,2188,-4574 $DEVICE_ID=1003
MM197 2 27 33 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-5122  $PIN_XY=2248,-5208,2218,-5122,2188,-5208 $DEVICE_ID=1003
MM198 2 28 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-5563  $PIN_XY=2248,-5498,2218,-5563,2188,-5498 $DEVICE_ID=1003
MM199 37 31 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-4660  $PIN_XY=2080,-4574,2050,-4660,2020,-4574 $DEVICE_ID=1003
MM200 33 31 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-5122  $PIN_XY=2080,-5208,2050,-5122,2020,-5208 $DEVICE_ID=1003
MM201 32 26 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-5563  $PIN_XY=2080,-5498,2050,-5563,2020,-5498 $DEVICE_ID=1003
MM202 2 30 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1378 $Y=-5202  $PIN_XY=1408,-5208,1378,-5202,1348,-5208 $DEVICE_ID=1003
MM203 28 30 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1210 $Y=-5202  $PIN_XY=1240,-5208,1210,-5202,1180,-5208 $DEVICE_ID=1003
MM204 2 34 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1042 $Y=-4681  $PIN_XY=1072,-4574,1042,-4681,1012,-4574 $DEVICE_ID=1003
MM205 2 30 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1042 $Y=-5101  $PIN_XY=1072,-5208,1042,-5101,1012,-5208 $DEVICE_ID=1003
MM206 30 34 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=874 $Y=-4681  $PIN_XY=904,-4574,874,-4681,844,-4574 $DEVICE_ID=1003
MM207 28 30 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=874 $Y=-5101  $PIN_XY=904,-5208,874,-5101,844,-5208 $DEVICE_ID=1003
XX30BB92C5772 16 17 35 31 66 73 inv $T=1324 716 1 0 $X=1324 $Y=126
XX30BB92C5773 15 14 29 26 65 75 inv $T=1324 1640 1 0 $X=1324 $Y=1050
XX30BB92C5774 16 14 36 27 66 75 inv $T=1324 590 0 0 $X=1324 $Y=590
XX30BB92C5775 8 2 19 41 37 76 62 69 nor $T=1872 -3902 1 0 $X=2500 $Y=-4494
XX30BB92C5776 13 6 21 43 39 77 64 71 nor $T=1872 -2054 1 0 $X=2500 $Y=-2646
XX30BB92C5777 5 7 20 42 38 78 61 70 nor $T=1872 -2978 1 0 $X=2500 $Y=-3570
XX30BB92C5778 3 2 18 33 32 79 60 68 nor $T=1872 -4826 1 0 $X=2500 $Y=-5418
XX30BB92C5779 10 12 22 47 40 80 63 72 nor $T=1872 -1130 1 0 $X=2500 $Y=-1722
XX30BB92C5780 11 9 23 48 44 81 67 74 nor $T=1872 -206 1 0 $X=2500 $Y=-798
XX30BB92C5781 15 14 25 50 46 82 65 75 nor $T=1872 1642 1 0 $X=2500 $Y=1050
XX30BB92C5782 16 17 24 49 45 83 66 73 nor $T=1872 718 1 0 $X=2500 $Y=126
XX30BB92C5783 5 6 39 31 28 92 61 71 nand $T=1410 -3334 0 0 $X=1827 $Y=-3106
XX30BB92C5784 13 6 43 29 36 93 64 71 nand $T=1410 -1828 1 0 $X=1827 $Y=-2646
XX30BB92C5785 5 7 42 31 36 94 61 70 nand $T=1410 -2752 1 0 $X=1827 $Y=-3570
XX30BB92C5786 8 7 38 26 28 95 62 70 nand $T=1410 -4258 0 0 $X=1827 $Y=-4030
XX30BB92C5787 4 2 32 26 28 112 59 68 nand $T=1410 -6106 0 0 $X=1827 $Y=-5878
XX30BB92C5788 3 2 37 31 28 96 60 69 nand $T=1410 -5182 0 0 $X=1827 $Y=-4954
XX30BB92C5789 8 2 41 29 27 97 62 69 nand $T=1410 -3676 1 0 $X=1827 $Y=-4494
XX30BB92C5790 3 2 33 31 27 98 60 68 nand $T=1410 -4600 1 0 $X=1827 $Y=-5418
XX30BB92C5791 11 17 45 35 28 99 67 73 nand $T=1410 -562 0 0 $X=1827 $Y=-334
XX30BB92C5792 13 12 40 35 28 100 64 72 nand $T=1410 -2410 0 0 $X=1827 $Y=-2182
XX30BB92C5793 10 12 47 26 27 101 63 72 nand $T=1410 -904 1 0 $X=1827 $Y=-1722
XX30BB92C5794 11 9 48 29 27 102 67 74 nand $T=1410 20 1 0 $X=1827 $Y=-798
XX30BB92C5795 10 9 44 35 28 103 63 74 nand $T=1410 -1486 0 0 $X=1827 $Y=-1258
XX30BB92C5796 16 17 49 26 36 104 66 73 nand $T=1410 944 1 0 $X=1827 $Y=126
XX30BB92C5797 15 14 50 29 36 105 65 75 nand $T=1410 1868 1 0 $X=1827 $Y=1050
XX30BB92C5798 16 14 46 35 28 106 66 75 nand $T=1410 362 0 0 $X=1827 $Y=590
XX30BB92C5799 6 5 51 84 21 39 61 71 buffer_highdrive $T=2498 -3104 0 0 $X=2500 $Y=-3106
XX30BB92C5800 2 3 52 85 19 37 60 69 buffer_highdrive $T=2498 -4952 0 0 $X=2500 $Y=-4954
XX30BB92C5801 12 13 53 86 22 40 64 72 buffer_highdrive $T=2498 -2180 0 0 $X=2500 $Y=-2182
XX30BB92C5802 9 10 54 87 23 44 63 74 buffer_highdrive $T=2498 -1256 0 0 $X=2500 $Y=-1258
XX30BB92C5803 2 4 55 88 18 32 59 68 buffer_highdrive $T=2498 -5876 0 0 $X=2500 $Y=-5878
XX30BB92C5804 7 8 56 89 20 38 62 70 buffer_highdrive $T=2498 -4028 0 0 $X=2500 $Y=-4030
XX30BB92C5805 14 16 57 90 25 46 66 75 buffer_highdrive $T=2498 592 0 0 $X=2500 $Y=590
XX30BB92C5806 17 11 58 91 24 45 67 73 buffer_highdrive $T=2498 -332 0 0 $X=2500 $Y=-334
XX30BB92C5807 3 2 28 30 60 68 invx4 $T=628 -4828 1 0 $X=652 $Y=-5418
XX30BB92C5808 3 2 30 34 60 69 invx4 $T=628 -4954 0 0 $X=652 $Y=-4954
XX30BB92C5809 15 14 _GENERATED_114 _GENERATED_113 65 75 sram_filler $T=1100 1640 0 180 $X=652 $Y=1050
XX30BB92C5810 16 14 _GENERATED_116 _GENERATED_115 66 75 sram_filler $T=648 590 0 0 $X=652 $Y=590
XX30BB92C5811 16 17 _GENERATED_118 _GENERATED_117 66 73 sram_filler $T=1100 716 0 180 $X=652 $Y=126
XX30BB92C5812 16 17 _GENERATED_120 _GENERATED_119 66 73 sram_filler $T=1436 716 0 180 $X=988 $Y=126
XX30BB92C5813 16 14 _GENERATED_122 _GENERATED_121 66 75 sram_filler $T=984 590 0 0 $X=988 $Y=590
XX30BB92C5814 15 14 _GENERATED_124 _GENERATED_123 65 75 sram_filler $T=1436 1640 0 180 $X=988 $Y=1050
XX30BB92C5815 4 2 _GENERATED_126 _GENERATED_125 59 68 sram_filler $T=648 -5878 0 0 $X=652 $Y=-5878
XX30BB92C5816 4 2 _GENERATED_128 _GENERATED_127 59 68 sram_filler $T=984 -5878 0 0 $X=988 $Y=-5878
XX30BB92C5817 4 2 _GENERATED_129 4 59 68 sram_filler $T=1320 -5878 0 0 $X=1324 $Y=-5878
XX30BB92C5818 4 2 2 _GENERATED_130 59 68 sram_filler $T=1488 -5878 0 0 $X=1492 $Y=-5878
XX30BB92C5819 11 17 _GENERATED_132 _GENERATED_131 67 73 sram_filler $T=648 -334 0 0 $X=652 $Y=-334
XX30BB92C5820 11 17 _GENERATED_134 _GENERATED_133 67 73 sram_filler $T=984 -334 0 0 $X=988 $Y=-334
XX30BB92C5821 11 17 _GENERATED_135 11 67 73 sram_filler $T=1320 -334 0 0 $X=1324 $Y=-334
XX30BB92C5822 11 17 17 _GENERATED_136 67 73 sram_filler $T=1488 -334 0 0 $X=1492 $Y=-334
XX30BB92C5823 10 9 _GENERATED_137 10 63 74 sram_filler $T=648 -1258 0 0 $X=652 $Y=-1258
XX30BB92C5824 10 9 9 _GENERATED_138 63 74 sram_filler $T=816 -1258 0 0 $X=820 $Y=-1258
XX30BB92C5825 10 9 _GENERATED_140 _GENERATED_139 63 74 sram_filler $T=1152 -1258 0 0 $X=1156 $Y=-1258
XX30BB92C5826 10 9 _GENERATED_142 _GENERATED_141 63 74 sram_filler $T=1488 -1258 0 0 $X=1492 $Y=-1258
XX30BB92C5827 11 9 9 _GENERATED_143 67 74 sram_filler $T=1100 -208 0 180 $X=652 $Y=-798
XX30BB92C5828 11 9 _GENERATED_144 11 67 74 sram_filler $T=1268 -208 0 180 $X=820 $Y=-798
XX30BB92C5829 11 9 _GENERATED_146 _GENERATED_145 67 74 sram_filler $T=1604 -208 0 180 $X=1156 $Y=-798
XX30BB92C5830 11 9 _GENERATED_148 _GENERATED_147 67 74 sram_filler $T=1940 -208 0 180 $X=1492 $Y=-798
XX30BB92C5831 10 12 _GENERATED_150 _GENERATED_149 63 72 sram_filler $T=1940 -1132 0 180 $X=1492 $Y=-1722
XX30BB92C5832 10 12 _GENERATED_152 _GENERATED_151 63 72 sram_filler $T=1604 -1132 0 180 $X=1156 $Y=-1722
XX30BB92C5833 10 12 _GENERATED_153 10 63 72 sram_filler $T=1268 -1132 0 180 $X=820 $Y=-1722
XX30BB92C5834 10 12 12 _GENERATED_154 63 72 sram_filler $T=1100 -1132 0 180 $X=652 $Y=-1722
XX30BB92C5835 13 12 _GENERATED_156 _GENERATED_155 64 72 sram_filler $T=1488 -2182 0 0 $X=1492 $Y=-2182
XX30BB92C5836 13 12 _GENERATED_158 _GENERATED_157 64 72 sram_filler $T=1152 -2182 0 0 $X=1156 $Y=-2182
XX30BB92C5837 13 12 12 _GENERATED_159 64 72 sram_filler $T=816 -2182 0 0 $X=820 $Y=-2182
XX30BB92C5838 13 12 _GENERATED_160 13 64 72 sram_filler $T=648 -2182 0 0 $X=652 $Y=-2182
XX30BB92C5839 13 6 6 _GENERATED_161 64 71 sram_filler $T=1100 -2056 0 180 $X=652 $Y=-2646
XX30BB92C5840 13 6 _GENERATED_162 13 64 71 sram_filler $T=1268 -2056 0 180 $X=820 $Y=-2646
XX30BB92C5841 13 6 _GENERATED_164 _GENERATED_163 64 71 sram_filler $T=1604 -2056 0 180 $X=1156 $Y=-2646
XX30BB92C5842 13 6 _GENERATED_166 _GENERATED_165 64 71 sram_filler $T=1940 -2056 0 180 $X=1492 $Y=-2646
XX30BB92C5843 5 6 _GENERATED_168 _GENERATED_167 61 71 sram_filler $T=648 -3106 0 0 $X=652 $Y=-3106
XX30BB92C5844 5 6 _GENERATED_170 _GENERATED_169 61 71 sram_filler $T=984 -3106 0 0 $X=988 $Y=-3106
XX30BB92C5845 5 6 _GENERATED_171 5 61 71 sram_filler $T=1320 -3106 0 0 $X=1324 $Y=-3106
XX30BB92C5846 5 6 6 _GENERATED_172 61 71 sram_filler $T=1488 -3106 0 0 $X=1492 $Y=-3106
XX30BB92C5847 5 7 _GENERATED_174 _GENERATED_173 61 70 sram_filler $T=1940 -2980 0 180 $X=1492 $Y=-3570
XX30BB92C5848 5 7 _GENERATED_176 _GENERATED_175 61 70 sram_filler $T=1604 -2980 0 180 $X=1156 $Y=-3570
XX30BB92C5849 5 7 _GENERATED_177 5 61 70 sram_filler $T=1268 -2980 0 180 $X=820 $Y=-3570
XX30BB92C5850 5 7 7 _GENERATED_178 61 70 sram_filler $T=1100 -2980 0 180 $X=652 $Y=-3570
XX30BB92C5851 8 7 7 _GENERATED_179 62 70 sram_filler $T=1488 -4030 0 0 $X=1492 $Y=-4030
XX30BB92C5852 8 7 _GENERATED_180 8 62 70 sram_filler $T=1320 -4030 0 0 $X=1324 $Y=-4030
XX30BB92C5853 8 7 _GENERATED_182 _GENERATED_181 62 70 sram_filler $T=984 -4030 0 0 $X=988 $Y=-4030
XX30BB92C5854 8 7 _GENERATED_184 _GENERATED_183 62 70 sram_filler $T=648 -4030 0 0 $X=652 $Y=-4030
XX30BB92C5855 8 2 2 _GENERATED_185 62 69 sram_filler $T=1100 -3904 0 180 $X=652 $Y=-4494
XX30BB92C5856 8 2 _GENERATED_186 8 62 69 sram_filler $T=1268 -3904 0 180 $X=820 $Y=-4494
XX30BB92C5857 8 2 _GENERATED_188 _GENERATED_187 62 69 sram_filler $T=1604 -3904 0 180 $X=1156 $Y=-4494
XX30BB92C5858 8 2 _GENERATED_190 _GENERATED_189 62 69 sram_filler $T=1940 -3904 0 180 $X=1492 $Y=-4494
XX30BB92C5859 13 6 _GENERATED_192 _GENERATED_191 64 71 sram_filler $T=3168 -2056 1 0 $X=3172 $Y=-2646
XX30BB92C5860 13 6 _GENERATED_194 _GENERATED_193 64 71 sram_filler $T=3840 -2056 1 0 $X=3844 $Y=-2646
XX30BB92C5861 13 6 _GENERATED_196 _GENERATED_195 64 71 sram_filler $T=3504 -2056 1 0 $X=3508 $Y=-2646
XX30BB92C5862 5 7 _GENERATED_198 _GENERATED_197 61 70 sram_filler $T=3840 -2980 1 0 $X=3844 $Y=-3570
XX30BB92C5863 5 7 _GENERATED_200 _GENERATED_199 61 70 sram_filler $T=3168 -2980 1 0 $X=3172 $Y=-3570
XX30BB92C5864 5 7 _GENERATED_202 _GENERATED_201 61 70 sram_filler $T=3504 -2980 1 0 $X=3508 $Y=-3570
XX30BB92C5865 8 2 _GENERATED_204 _GENERATED_203 62 69 sram_filler $T=3168 -3904 1 0 $X=3172 $Y=-4494
XX30BB92C5866 8 2 _GENERATED_206 _GENERATED_205 62 69 sram_filler $T=3840 -3904 1 0 $X=3844 $Y=-4494
XX30BB92C5867 8 2 _GENERATED_208 _GENERATED_207 62 69 sram_filler $T=3504 -3904 1 0 $X=3508 $Y=-4494
XX30BB92C5868 3 2 _GENERATED_210 _GENERATED_209 60 68 sram_filler $T=3840 -4828 1 0 $X=3844 $Y=-5418
XX30BB92C5869 3 2 _GENERATED_212 _GENERATED_211 60 68 sram_filler $T=3168 -4828 1 0 $X=3172 $Y=-5418
XX30BB92C5870 3 2 _GENERATED_214 _GENERATED_213 60 68 sram_filler $T=3504 -4828 1 0 $X=3508 $Y=-5418
XX30BB92C5871 10 12 _GENERATED_216 _GENERATED_215 63 72 sram_filler $T=3504 -1132 1 0 $X=3508 $Y=-1722
XX30BB92C5872 10 12 _GENERATED_218 _GENERATED_217 63 72 sram_filler $T=3168 -1132 1 0 $X=3172 $Y=-1722
XX30BB92C5873 10 12 _GENERATED_220 _GENERATED_219 63 72 sram_filler $T=3840 -1132 1 0 $X=3844 $Y=-1722
XX30BB92C5874 11 9 _GENERATED_222 _GENERATED_221 67 74 sram_filler $T=3504 -208 1 0 $X=3508 $Y=-798
XX30BB92C5875 11 9 _GENERATED_224 _GENERATED_223 67 74 sram_filler $T=3840 -208 1 0 $X=3844 $Y=-798
XX30BB92C5876 11 9 _GENERATED_226 _GENERATED_225 67 74 sram_filler $T=3168 -208 1 0 $X=3172 $Y=-798
XX30BB92C5877 16 17 _GENERATED_228 _GENERATED_227 66 73 sram_filler $T=3168 716 1 0 $X=3172 $Y=126
XX30BB92C5878 16 17 _GENERATED_230 _GENERATED_229 66 73 sram_filler $T=3840 716 1 0 $X=3844 $Y=126
XX30BB92C5879 15 14 _GENERATED_232 _GENERATED_231 65 75 sram_filler $T=3840 1640 1 0 $X=3844 $Y=1050
XX30BB92C5880 15 14 _GENERATED_234 _GENERATED_233 65 75 sram_filler $T=3168 1640 1 0 $X=3172 $Y=1050
XX30BB92C5881 15 14 _GENERATED_236 _GENERATED_235 65 75 sram_filler $T=3504 1640 1 0 $X=3508 $Y=1050
XX30BB92C5882 16 17 _GENERATED_238 _GENERATED_237 66 73 sram_filler $T=3504 716 1 0 $X=3508 $Y=126
XX30BB92C5883 3 2 _GENERATED_240 _GENERATED_239 60 68 sram_filler $T=1488 -4828 1 0 $X=1492 $Y=-5418
XX30BB92C5884 3 2 _GENERATED_242 _GENERATED_241 60 69 sram_filler $T=1488 -4954 0 0 $X=1492 $Y=-4954
.ends static_row_decoder_3by8
.subckt WLRef_PC 2 3 4 5 6 7 8 9 10 12 15
+	19 22 24 26 27 29 33 34 36 37 38
+	42 49 50 51 58 59 60 61 62 63 64
+	71
*.floating_nets 70
MM1 8 35 40 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5770 $Y=1241  $PIN_XY=5800,1136,5770,1241,5740,1136 $DEVICE_ID=1001
MM2 34 41 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5602 $Y=1661  $PIN_XY=5632,1766,5602,1661,5572,1766 $DEVICE_ID=1001
MM3 35 39 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5602 $Y=737  $PIN_XY=5632,842,5602,737,5572,842 $DEVICE_ID=1001
MM4 8 40 32 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5266 $Y=1241  $PIN_XY=5296,1136,5266,1241,5236,1136 $DEVICE_ID=1001
MM5 41 32 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5098 $Y=1661  $PIN_XY=5128,1766,5098,1661,5068,1766 $DEVICE_ID=1001
MM6 39 30 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5098 $Y=737  $PIN_XY=5128,842,5098,737,5068,842 $DEVICE_ID=1001
MM7 8 31 44 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4762 $Y=1241  $PIN_XY=4792,1136,4762,1241,4732,1136 $DEVICE_ID=1001
MM8 31 45 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4594 $Y=1682  $PIN_XY=4624,1766,4594,1682,4564,1766 $DEVICE_ID=1001
MM9 30 43 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4594 $Y=737  $PIN_XY=4624,842,4594,737,4564,842 $DEVICE_ID=1001
MM10 2 23 38 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4426 $Y=2165  $PIN_XY=4456,2060,4426,2165,4396,2060 $DEVICE_ID=1001
MM11 38 23 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4258 $Y=2165  $PIN_XY=4288,2060,4258,2165,4228,2060 $DEVICE_ID=1001
MM12 8 44 28 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4258 $Y=1241  $PIN_XY=4288,1136,4258,1241,4228,1136 $DEVICE_ID=1001
MM13 45 22 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4090 $Y=1661  $PIN_XY=4120,1766,4090,1661,4060,1766 $DEVICE_ID=1001
MM14 43 28 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4090 $Y=737  $PIN_XY=4120,842,4090,737,4060,842 $DEVICE_ID=1001
MM15 2 12 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3754 $Y=2144  $PIN_XY=3784,2060,3754,2144,3724,2060 $DEVICE_ID=1001
MM16 2 24 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3754 $Y=1703  $PIN_XY=3784,1766,3754,1703,3724,1766 $DEVICE_ID=1001
MM17 23 25 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3586 $Y=2165  $PIN_XY=3616,2060,3586,2165,3556,2060 $DEVICE_ID=1001
MM18 2 21 48 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3250 $Y=1661  $PIN_XY=3280,1766,3250,1661,3220,1766 $DEVICE_ID=1001
MM19 8 20 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3250 $Y=737  $PIN_XY=3280,842,3250,737,3220,842 $DEVICE_ID=1001
MM20 21 67 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3082 $Y=2144  $PIN_XY=3112,2060,3082,2144,3052,2060 $DEVICE_ID=1001
MM21 20 54 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3082 $Y=1241  $PIN_XY=3112,1136,3082,1241,3052,1136 $DEVICE_ID=1001
MM22 2 48 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2746 $Y=1661  $PIN_XY=2776,1766,2746,1661,2716,1766 $DEVICE_ID=1001
MM23 8 55 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2746 $Y=737  $PIN_XY=2776,842,2746,737,2716,842 $DEVICE_ID=1001
MM24 67 17 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2578 $Y=2144  $PIN_XY=2608,2060,2578,2144,2548,2060 $DEVICE_ID=1001
MM25 54 16 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2578 $Y=1241  $PIN_XY=2608,1136,2578,1241,2548,1136 $DEVICE_ID=1001
MM26 2 19 47 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2242 $Y=1661  $PIN_XY=2272,1766,2242,1661,2212,1766 $DEVICE_ID=1001
MM27 8 18 56 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2242 $Y=737  $PIN_XY=2272,842,2242,737,2212,842 $DEVICE_ID=1001
MM28 17 68 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2074 $Y=2144  $PIN_XY=2104,2060,2074,2144,2044,2060 $DEVICE_ID=1001
MM29 16 53 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2074 $Y=1241  $PIN_XY=2104,1136,2074,1241,2044,1136 $DEVICE_ID=1001
MM30 2 47 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1738 $Y=1661  $PIN_XY=1768,1766,1738,1661,1708,1766 $DEVICE_ID=1001
MM31 8 56 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1738 $Y=737  $PIN_XY=1768,842,1738,737,1708,842 $DEVICE_ID=1001
MM32 68 12 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1570 $Y=2144  $PIN_XY=1600,2060,1570,2144,1540,2060 $DEVICE_ID=1001
MM33 53 11 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1570 $Y=1241  $PIN_XY=1600,1136,1570,1241,1540,1136 $DEVICE_ID=1001
MM34 2 14 46 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1234 $Y=1661  $PIN_XY=1264,1766,1234,1661,1204,1766 $DEVICE_ID=1001
MM35 8 13 57 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1234 $Y=737  $PIN_XY=1264,842,1234,737,1204,842 $DEVICE_ID=1001
MM36 12 69 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1066 $Y=2144  $PIN_XY=1096,2060,1066,2144,1036,2060 $DEVICE_ID=1001
MM37 11 52 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1066 $Y=1241  $PIN_XY=1096,1136,1066,1241,1036,1136 $DEVICE_ID=1001
MM38 2 46 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=730 $Y=1661  $PIN_XY=760,1766,730,1661,700,1766 $DEVICE_ID=1001
MM39 8 57 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=730 $Y=737  $PIN_XY=760,842,730,737,700,842 $DEVICE_ID=1001
MM40 69 24 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=562 $Y=2144  $PIN_XY=592,2060,562,2144,532,2060 $DEVICE_ID=1001
MM41 52 25 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=562 $Y=1241  $PIN_XY=592,1136,562,1241,532,1136 $DEVICE_ID=1001
MM42 3 41 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5770 $Y=1581  $PIN_XY=5800,1596,5770,1581,5740,1596 $DEVICE_ID=1003
MM43 3 35 40 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5770 $Y=1241  $PIN_XY=5800,1306,5770,1241,5740,1306 $DEVICE_ID=1003
MM44 5 39 35 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5770 $Y=678  $PIN_XY=5800,672,5770,678,5740,672 $DEVICE_ID=1003
MM45 34 41 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5602 $Y=1661  $PIN_XY=5632,1596,5602,1661,5572,1596 $DEVICE_ID=1003
MM46 40 35 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5602 $Y=1321  $PIN_XY=5632,1306,5602,1321,5572,1306 $DEVICE_ID=1003
MM47 35 39 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5602 $Y=737  $PIN_XY=5632,672,5602,737,5572,672 $DEVICE_ID=1003
MM48 33 22 65 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5602 $Y=317  $PIN_XY=5632,382,5602,317,5572,382 $DEVICE_ID=1003
MM49 65 34 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5434 $Y=296  $PIN_XY=5464,382,5434,296,5404,382 $DEVICE_ID=1003
MM50 3 32 41 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5266 $Y=1581  $PIN_XY=5296,1596,5266,1581,5236,1596 $DEVICE_ID=1003
MM51 3 40 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5266 $Y=1241  $PIN_XY=5296,1306,5266,1241,5236,1306 $DEVICE_ID=1003
MM52 5 30 39 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5266 $Y=678  $PIN_XY=5296,672,5266,678,5236,672 $DEVICE_ID=1003
MM53 41 32 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5098 $Y=1661  $PIN_XY=5128,1596,5098,1661,5068,1596 $DEVICE_ID=1003
MM54 32 40 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5098 $Y=1321  $PIN_XY=5128,1306,5098,1321,5068,1306 $DEVICE_ID=1003
MM55 39 30 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5098 $Y=737  $PIN_XY=5128,672,5098,737,5068,672 $DEVICE_ID=1003
MM56 5 33 37 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5098 $Y=397  $PIN_XY=5128,382,5098,397,5068,382 $DEVICE_ID=1003
MM57 37 33 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4930 $Y=376  $PIN_XY=4960,382,4930,376,4900,382 $DEVICE_ID=1003
MM58 6 27 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=2585  $PIN_XY=4792,2520,4762,2585,4732,2520 $DEVICE_ID=1003
MM59 6 23 38 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=2245  $PIN_XY=4792,2230,4762,2245,4732,2230 $DEVICE_ID=1003
MM60 3 45 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=1581  $PIN_XY=4792,1596,4762,1581,4732,1596 $DEVICE_ID=1003
MM61 3 31 44 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=1241  $PIN_XY=4792,1306,4762,1241,4732,1306 $DEVICE_ID=1003
MM62 5 43 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=657  $PIN_XY=4792,672,4762,657,4732,672 $DEVICE_ID=1003
MM63 5 33 37 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4762 $Y=317  $PIN_XY=4792,382,4762,317,4732,382 $DEVICE_ID=1003
MM64 36 27 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4594 $Y=2585  $PIN_XY=4624,2520,4594,2585,4564,2520 $DEVICE_ID=1003
MM65 38 23 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4594 $Y=2245  $PIN_XY=4624,2230,4594,2245,4564,2230 $DEVICE_ID=1003
MM66 31 45 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4594 $Y=1682  $PIN_XY=4624,1596,4594,1682,4564,1596 $DEVICE_ID=1003
MM67 44 31 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4594 $Y=1321  $PIN_XY=4624,1306,4594,1321,4564,1306 $DEVICE_ID=1003
MM68 30 43 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4594 $Y=737  $PIN_XY=4624,672,4594,737,4564,672 $DEVICE_ID=1003
MM69 37 33 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4594 $Y=317  $PIN_XY=4624,382,4594,317,4564,382 $DEVICE_ID=1003
MM70 6 27 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4426 $Y=2505  $PIN_XY=4456,2520,4426,2505,4396,2520 $DEVICE_ID=1003
MM71 6 23 38 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4426 $Y=2165  $PIN_XY=4456,2230,4426,2165,4396,2230 $DEVICE_ID=1003
MM72 36 27 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4258 $Y=2505  $PIN_XY=4288,2520,4258,2505,4228,2520 $DEVICE_ID=1003
MM73 38 23 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4258 $Y=2165  $PIN_XY=4288,2230,4258,2165,4228,2230 $DEVICE_ID=1003
MM74 3 22 45 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4258 $Y=1581  $PIN_XY=4288,1596,4258,1581,4228,1596 $DEVICE_ID=1003
MM75 3 44 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4258 $Y=1241  $PIN_XY=4288,1306,4258,1241,4228,1306 $DEVICE_ID=1003
MM76 5 28 43 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4258 $Y=657  $PIN_XY=4288,672,4258,657,4228,672 $DEVICE_ID=1003
MM77 5 42 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4258 $Y=397  $PIN_XY=4288,382,4258,397,4228,382 $DEVICE_ID=1003
MM78 45 22 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4090 $Y=1661  $PIN_XY=4120,1596,4090,1661,4060,1596 $DEVICE_ID=1003
MM79 28 44 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4090 $Y=1321  $PIN_XY=4120,1306,4090,1321,4060,1306 $DEVICE_ID=1003
MM80 43 28 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4090 $Y=737  $PIN_XY=4120,672,4090,737,4060,672 $DEVICE_ID=1003
MM81 29 42 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4090 $Y=317  $PIN_XY=4120,382,4090,317,4060,382 $DEVICE_ID=1003
MM82 6 19 27 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3754 $Y=2585  $PIN_XY=3784,2520,3754,2585,3724,2520 $DEVICE_ID=1003
MM83 23 12 66 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3754 $Y=2144  $PIN_XY=3784,2230,3754,2144,3724,2230 $DEVICE_ID=1003
MM84 3 24 22 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3754 $Y=1703  $PIN_XY=3784,1596,3754,1703,3724,1596 $DEVICE_ID=1003
MM85 5 26 42 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3754 $Y=376  $PIN_XY=3784,382,3754,376,3724,382 $DEVICE_ID=1003
MM86 27 12 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3586 $Y=2585  $PIN_XY=3616,2520,3586,2585,3556,2520 $DEVICE_ID=1003
MM87 66 25 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3586 $Y=2165  $PIN_XY=3616,2230,3586,2165,3556,2230 $DEVICE_ID=1003
MM88 22 24 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3586 $Y=1602  $PIN_XY=3616,1596,3586,1602,3556,1596 $DEVICE_ID=1003
MM89 42 26 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3586 $Y=296  $PIN_XY=3616,382,3586,296,3556,382 $DEVICE_ID=1003
MM90 6 67 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3250 $Y=2224  $PIN_XY=3280,2230,3250,2224,3220,2230 $DEVICE_ID=1003
MM91 3 21 48 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3250 $Y=1661  $PIN_XY=3280,1596,3250,1661,3220,1596 $DEVICE_ID=1003
MM92 3 54 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3250 $Y=1321  $PIN_XY=3280,1306,3250,1321,3220,1306 $DEVICE_ID=1003
MM93 5 20 55 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3250 $Y=737  $PIN_XY=3280,672,3250,737,3220,672 $DEVICE_ID=1003
MM94 5 51 26 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3250 $Y=397  $PIN_XY=3280,382,3250,397,3220,382 $DEVICE_ID=1003
MM95 21 67 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3082 $Y=2144  $PIN_XY=3112,2230,3082,2144,3052,2230 $DEVICE_ID=1003
MM96 48 21 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3082 $Y=1581  $PIN_XY=3112,1596,3082,1581,3052,1596 $DEVICE_ID=1003
MM97 20 54 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3082 $Y=1241  $PIN_XY=3112,1306,3082,1241,3052,1306 $DEVICE_ID=1003
MM98 55 20 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3082 $Y=657  $PIN_XY=3112,672,3082,657,3052,672 $DEVICE_ID=1003
MM99 26 51 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3082 $Y=317  $PIN_XY=3112,382,3082,317,3052,382 $DEVICE_ID=1003
MM100 6 17 67 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2746 $Y=2224  $PIN_XY=2776,2230,2746,2224,2716,2230 $DEVICE_ID=1003
MM101 3 48 19 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2746 $Y=1661  $PIN_XY=2776,1596,2746,1661,2716,1596 $DEVICE_ID=1003
MM102 3 16 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2746 $Y=1321  $PIN_XY=2776,1306,2746,1321,2716,1306 $DEVICE_ID=1003
MM103 5 55 18 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2746 $Y=737  $PIN_XY=2776,672,2746,737,2716,672 $DEVICE_ID=1003
MM104 5 15 51 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2746 $Y=397  $PIN_XY=2776,382,2746,397,2716,382 $DEVICE_ID=1003
MM105 67 17 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2578 $Y=2144  $PIN_XY=2608,2230,2578,2144,2548,2230 $DEVICE_ID=1003
MM106 19 48 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2578 $Y=1581  $PIN_XY=2608,1596,2578,1581,2548,1596 $DEVICE_ID=1003
MM107 54 16 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2578 $Y=1241  $PIN_XY=2608,1306,2578,1241,2548,1306 $DEVICE_ID=1003
MM108 18 55 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2578 $Y=657  $PIN_XY=2608,672,2578,657,2548,672 $DEVICE_ID=1003
MM109 51 15 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2578 $Y=317  $PIN_XY=2608,382,2578,317,2548,382 $DEVICE_ID=1003
MM110 6 68 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2242 $Y=2224  $PIN_XY=2272,2230,2242,2224,2212,2230 $DEVICE_ID=1003
MM111 3 19 47 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2242 $Y=1661  $PIN_XY=2272,1596,2242,1661,2212,1596 $DEVICE_ID=1003
MM112 3 53 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2242 $Y=1321  $PIN_XY=2272,1306,2242,1321,2212,1306 $DEVICE_ID=1003
MM113 5 18 56 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2242 $Y=737  $PIN_XY=2272,672,2242,737,2212,672 $DEVICE_ID=1003
MM114 5 50 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2242 $Y=397  $PIN_XY=2272,382,2242,397,2212,382 $DEVICE_ID=1003
MM115 17 68 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2074 $Y=2144  $PIN_XY=2104,2230,2074,2144,2044,2230 $DEVICE_ID=1003
MM116 47 19 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2074 $Y=1581  $PIN_XY=2104,1596,2074,1581,2044,1596 $DEVICE_ID=1003
MM117 16 53 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2074 $Y=1241  $PIN_XY=2104,1306,2074,1241,2044,1306 $DEVICE_ID=1003
MM118 56 18 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2074 $Y=657  $PIN_XY=2104,672,2074,657,2044,672 $DEVICE_ID=1003
MM119 15 50 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2074 $Y=317  $PIN_XY=2104,382,2074,317,2044,382 $DEVICE_ID=1003
MM120 6 12 68 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1738 $Y=2224  $PIN_XY=1768,2230,1738,2224,1708,2230 $DEVICE_ID=1003
MM121 3 47 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1738 $Y=1661  $PIN_XY=1768,1596,1738,1661,1708,1596 $DEVICE_ID=1003
MM122 3 11 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1738 $Y=1321  $PIN_XY=1768,1306,1738,1321,1708,1306 $DEVICE_ID=1003
MM123 5 56 13 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1738 $Y=737  $PIN_XY=1768,672,1738,737,1708,672 $DEVICE_ID=1003
MM124 5 10 50 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1738 $Y=397  $PIN_XY=1768,382,1738,397,1708,382 $DEVICE_ID=1003
MM125 68 12 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1570 $Y=2144  $PIN_XY=1600,2230,1570,2144,1540,2230 $DEVICE_ID=1003
MM126 14 47 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1570 $Y=1581  $PIN_XY=1600,1596,1570,1581,1540,1596 $DEVICE_ID=1003
MM127 53 11 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1570 $Y=1241  $PIN_XY=1600,1306,1570,1241,1540,1306 $DEVICE_ID=1003
MM128 13 56 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1570 $Y=657  $PIN_XY=1600,672,1570,657,1540,672 $DEVICE_ID=1003
MM129 50 10 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1570 $Y=317  $PIN_XY=1600,382,1570,317,1540,382 $DEVICE_ID=1003
MM130 6 69 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1234 $Y=2224  $PIN_XY=1264,2230,1234,2224,1204,2230 $DEVICE_ID=1003
MM131 3 14 46 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1234 $Y=1661  $PIN_XY=1264,1596,1234,1661,1204,1596 $DEVICE_ID=1003
MM132 3 52 11 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1234 $Y=1321  $PIN_XY=1264,1306,1234,1321,1204,1306 $DEVICE_ID=1003
MM133 5 13 57 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1234 $Y=737  $PIN_XY=1264,672,1234,737,1204,672 $DEVICE_ID=1003
MM134 5 49 10 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1234 $Y=397  $PIN_XY=1264,382,1234,397,1204,382 $DEVICE_ID=1003
MM135 12 69 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1066 $Y=2144  $PIN_XY=1096,2230,1066,2144,1036,2230 $DEVICE_ID=1003
MM136 46 14 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1066 $Y=1581  $PIN_XY=1096,1596,1066,1581,1036,1596 $DEVICE_ID=1003
MM137 11 52 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1066 $Y=1241  $PIN_XY=1096,1306,1066,1241,1036,1306 $DEVICE_ID=1003
MM138 57 13 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1066 $Y=657  $PIN_XY=1096,672,1066,657,1036,672 $DEVICE_ID=1003
MM139 10 49 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1066 $Y=317  $PIN_XY=1096,382,1066,317,1036,382 $DEVICE_ID=1003
MM140 6 24 69 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=730 $Y=2224  $PIN_XY=760,2230,730,2224,700,2230 $DEVICE_ID=1003
MM141 3 46 25 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=730 $Y=1661  $PIN_XY=760,1596,730,1661,700,1596 $DEVICE_ID=1003
MM142 3 25 52 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=730 $Y=1321  $PIN_XY=760,1306,730,1321,700,1306 $DEVICE_ID=1003
MM143 5 57 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=730 $Y=737  $PIN_XY=760,672,730,737,700,672 $DEVICE_ID=1003
MM144 5 9 49 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=730 $Y=397  $PIN_XY=760,382,730,397,700,382 $DEVICE_ID=1003
MM145 69 24 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=562 $Y=2144  $PIN_XY=592,2230,562,2144,532,2230 $DEVICE_ID=1003
MM146 25 46 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=562 $Y=1581  $PIN_XY=592,1596,562,1581,532,1596 $DEVICE_ID=1003
MM147 52 25 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=562 $Y=1241  $PIN_XY=592,1306,562,1241,532,1306 $DEVICE_ID=1003
MM148 9 57 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=562 $Y=657  $PIN_XY=592,672,562,657,532,672 $DEVICE_ID=1003
MM149 49 9 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=562 $Y=317  $PIN_XY=592,382,562,317,532,382 $DEVICE_ID=1003
XX30BB92C5885 2 3 22 24 59 62 inv $T=3976 1976 0 180 $X=3364 $Y=1386
XX30BB92C5886 4 5 33 22 34 65 61 63 nor $T=4584 0 0 0 $X=5212 $Y=2
XX30BB92C5887 2 6 23 12 25 66 59 64 nor $T=2736 1848 0 0 $X=3364 $Y=1850
XX30BB92C5888 7 6 27 12 19 71 58 64 nand $T=2946 3128 1 0 $X=3364 $Y=2310
XX30BB92C5889 7 6 36 27 58 64 invx4 $T=5008 2900 0 180 $X=4035 $Y=2310
XX30BB92C5890 4 5 37 33 61 63 invx4 $T=4348 2 0 0 $X=4372 $Y=2
XX30BB92C5891 2 6 38 23 59 64 invx4 $T=4012 1850 0 0 $X=4036 $Y=1850
XX30BB92C5892 8 5 39 35 30 60 63 buffer $T=4796 1054 1 0 $X=4876 $Y=462
XX30BB92C5893 8 3 40 32 35 60 62 buffer $T=6072 924 1 180 $X=4876 $Y=926
XX30BB92C5894 2 3 41 34 32 59 62 buffer $T=4796 1978 1 0 $X=4876 $Y=1386
XX30BB92C5895 4 5 42 29 26 61 63 buffer $T=3284 0 0 0 $X=3364 $Y=2
XX30BB92C5896 8 5 43 30 28 60 63 buffer $T=3788 1054 1 0 $X=3868 $Y=462
XX30BB92C5897 8 3 44 28 31 60 62 buffer $T=5064 924 1 180 $X=3868 $Y=926
XX30BB92C5898 2 3 45 31 22 59 62 buffer $T=3788 1978 1 0 $X=3868 $Y=1386
XX30BB92C5899 2 3 46 25 14 59 62 buffer $T=1536 1978 0 180 $X=340 $Y=1386
XX30BB92C5900 2 3 47 14 19 59 62 buffer $T=2544 1978 0 180 $X=1348 $Y=1386
XX30BB92C5901 2 3 48 19 21 59 62 buffer $T=3552 1978 0 180 $X=2356 $Y=1386
XX30BB92C5902 2 6 67 21 17 59 64 buffer $T=2276 1848 0 0 $X=2356 $Y=1850
XX30BB92C5903 2 6 68 17 12 59 64 buffer $T=1268 1848 0 0 $X=1348 $Y=1850
XX30BB92C5904 2 6 69 12 24 59 64 buffer $T=260 1848 0 0 $X=340 $Y=1850
XX30BB92C5905 4 5 49 10 9 61 63 buffer $T=260 0 0 0 $X=340 $Y=2
XX30BB92C5906 4 5 50 15 10 61 63 buffer $T=1268 0 0 0 $X=1348 $Y=2
XX30BB92C5907 4 5 51 26 15 61 63 buffer $T=2276 0 0 0 $X=2356 $Y=2
XX30BB92C5908 8 3 52 11 25 60 62 buffer $T=260 924 0 0 $X=340 $Y=926
XX30BB92C5909 8 3 53 16 11 60 62 buffer $T=1268 924 0 0 $X=1348 $Y=926
XX30BB92C5910 8 3 54 20 16 60 62 buffer $T=2276 924 0 0 $X=2356 $Y=926
XX30BB92C5911 8 5 55 18 20 60 63 buffer $T=3552 1054 0 180 $X=2356 $Y=462
XX30BB92C5912 8 5 56 13 18 60 63 buffer $T=2544 1054 0 180 $X=1348 $Y=462
XX30BB92C5913 8 5 57 9 13 60 63 buffer $T=1536 1054 0 180 $X=340 $Y=462
XX30BB92C5914 7 6 _GENERATED_73 _GENERATED_72 58 64 sram_filler $T=788 2900 0 180 $X=340 $Y=2310
XX30BB92C5915 7 6 _GENERATED_75 _GENERATED_74 58 64 sram_filler $T=1124 2900 0 180 $X=676 $Y=2310
XX30BB92C5916 7 6 _GENERATED_77 _GENERATED_76 58 64 sram_filler $T=1460 2900 0 180 $X=1012 $Y=2310
XX30BB92C5917 7 6 _GENERATED_79 _GENERATED_78 58 64 sram_filler $T=1796 2900 0 180 $X=1348 $Y=2310
XX30BB92C5918 7 6 _GENERATED_81 _GENERATED_80 58 64 sram_filler $T=2132 2900 0 180 $X=1684 $Y=2310
XX30BB92C5919 7 6 _GENERATED_83 _GENERATED_82 58 64 sram_filler $T=2468 2900 0 180 $X=2020 $Y=2310
XX30BB92C5920 7 6 _GENERATED_85 _GENERATED_84 58 64 sram_filler $T=2804 2900 0 180 $X=2356 $Y=2310
XX30BB92C5921 7 6 _GENERATED_87 _GENERATED_86 58 64 sram_filler $T=3140 2900 0 180 $X=2692 $Y=2310
XX30BB92C5922 7 6 _GENERATED_89 _GENERATED_88 58 64 sram_filler $T=3476 2900 0 180 $X=3028 $Y=2310
XX30BB92C5923 7 6 _GENERATED_91 _GENERATED_90 58 64 sram_filler $T=5996 2900 0 180 $X=5548 $Y=2310
XX30BB92C5924 7 6 _GENERATED_93 _GENERATED_92 58 64 sram_filler $T=5660 2900 0 180 $X=5212 $Y=2310
XX30BB92C5925 7 6 _GENERATED_95 _GENERATED_94 58 64 sram_filler $T=5324 2900 0 180 $X=4875 $Y=2310
XX30BB92C5926 2 6 _GENERATED_97 _GENERATED_96 59 64 sram_filler $T=5544 1850 0 0 $X=5548 $Y=1850
XX30BB92C5927 2 6 _GENERATED_99 _GENERATED_98 59 64 sram_filler $T=5208 1850 0 0 $X=5212 $Y=1850
XX30BB92C5928 2 6 _GENERATED_101 _GENERATED_100 59 64 sram_filler $T=4872 1850 0 0 $X=4875 $Y=1850
XX30BB92C5929 8 5 5 _GENERATED_102 60 63 sram_filler $T=3812 1052 0 180 $X=3364 $Y=462
XX30BB92C5930 8 5 _GENERATED_103 8 60 63 sram_filler $T=3980 1052 0 180 $X=3532 $Y=462
XX30BB92C5931 8 3 3 _GENERATED_104 60 62 sram_filler $T=3528 926 0 0 $X=3532 $Y=926
XX30BB92C5932 8 3 _GENERATED_105 8 60 62 sram_filler $T=3360 926 0 0 $X=3364 $Y=926
.ends WLRef_PC
.subckt agen_unit 2 3 4 5 6 7 8 9 10 14 15
+	18 19 20 23 26 27 28 29 30 31 32
+	33 35 37 38 39 40 41 42 43 44 45
+	46 47 59 60 61
MM1 8 23 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=1895  $PIN_XY=3782,1832,3752,1895,3722,1832 $DEVICE_ID=1001
MM2 8 25 26 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=1454  $PIN_XY=3782,1538,3752,1454,3722,1538 $DEVICE_ID=1001
MM3 10 21 32 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=992  $PIN_XY=3782,908,3752,992,3722,908 $DEVICE_ID=1001
MM4 10 36 31 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=530  $PIN_XY=3782,614,3752,530,3722,614 $DEVICE_ID=1001
MM5 3 24 30 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=68  $PIN_XY=3782,-16,3752,68,3722,-16 $DEVICE_ID=1001
MM6 3 22 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=-394  $PIN_XY=3782,-310,3752,-394,3722,-310 $DEVICE_ID=1001
MM7 5 34 28 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=-856  $PIN_XY=3782,-940,3752,-856,3722,-940 $DEVICE_ID=1001
MM8 5 35 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=-1297  $PIN_XY=3782,-1234,3752,-1297,3722,-1234 $DEVICE_ID=1001
MM9 33 23 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=1895  $PIN_XY=3614,1832,3584,1895,3554,1832 $DEVICE_ID=1001
MM10 26 25 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=1454  $PIN_XY=3614,1538,3584,1454,3554,1538 $DEVICE_ID=1001
MM11 32 21 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=992  $PIN_XY=3614,908,3584,992,3554,908 $DEVICE_ID=1001
MM12 31 36 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=530  $PIN_XY=3614,614,3584,530,3554,614 $DEVICE_ID=1001
MM13 30 24 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=68  $PIN_XY=3614,-16,3584,68,3554,-16 $DEVICE_ID=1001
MM14 29 22 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-394  $PIN_XY=3614,-310,3584,-394,3554,-310 $DEVICE_ID=1001
MM15 28 34 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-856  $PIN_XY=3614,-940,3584,-856,3554,-940 $DEVICE_ID=1001
MM16 27 35 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-1297  $PIN_XY=3614,-1234,3584,-1297,3554,-1234 $DEVICE_ID=1001
MM17 10 12 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=971  $PIN_XY=3278,908,3248,971,3218,908 $DEVICE_ID=1001
MM18 10 17 36 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=551  $PIN_XY=3278,614,3248,551,3218,614 $DEVICE_ID=1001
MM19 5 11 34 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=-877  $PIN_XY=3278,-940,3248,-877,3218,-940 $DEVICE_ID=1001
MM20 5 15 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=-1297  $PIN_XY=3278,-1234,3248,-1297,3218,-1234 $DEVICE_ID=1001
MM21 23 20 58 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=1895  $PIN_XY=3110,1832,3080,1895,3050,1832 $DEVICE_ID=1001
MM22 25 20 57 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=1454  $PIN_XY=3110,1538,3080,1454,3050,1538 $DEVICE_ID=1001
MM23 21 20 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=992  $PIN_XY=3110,908,3080,992,3050,908 $DEVICE_ID=1001
MM24 36 20 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=530  $PIN_XY=3110,614,3080,530,3050,614 $DEVICE_ID=1001
MM25 24 20 56 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=68  $PIN_XY=3110,-16,3080,68,3050,-16 $DEVICE_ID=1001
MM26 22 20 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=-394  $PIN_XY=3110,-310,3080,-394,3050,-310 $DEVICE_ID=1001
MM27 34 20 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=-856  $PIN_XY=3110,-940,3080,-856,3050,-940 $DEVICE_ID=1001
MM28 35 20 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=-1297  $PIN_XY=3110,-1234,3080,-1297,3050,-1234 $DEVICE_ID=1001
MM29 58 18 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=1895  $PIN_XY=2942,1832,2912,1895,2882,1832 $DEVICE_ID=1001
MM30 57 14 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=1475  $PIN_XY=2942,1538,2912,1475,2882,1538 $DEVICE_ID=1001
MM31 56 16 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=47  $PIN_XY=2942,-16,2912,47,2882,-16 $DEVICE_ID=1001
MM32 55 13 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=-373  $PIN_XY=2942,-310,2912,-373,2882,-310 $DEVICE_ID=1001
MM33 20 19 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2408 $Y=992  $PIN_XY=2438,908,2408,992,2378,908 $DEVICE_ID=1001
MM34 8 12 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2072 $Y=1454  $PIN_XY=2102,1538,2072,1454,2042,1538 $DEVICE_ID=1001
MM35 3 11 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2072 $Y=-394  $PIN_XY=2102,-310,2072,-394,2042,-310 $DEVICE_ID=1001
MM36 18 14 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1904 $Y=1916  $PIN_XY=1934,1832,1904,1916,1874,1832 $DEVICE_ID=1001
MM37 16 13 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1904 $Y=68  $PIN_XY=1934,-16,1904,68,1874,-16 $DEVICE_ID=1001
MM38 7 25 26 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=1353  $PIN_XY=4118,1368,4088,1353,4058,1368 $DEVICE_ID=1003
MM39 7 21 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=1093  $PIN_XY=4118,1078,4088,1093,4058,1078 $DEVICE_ID=1003
MM40 4 36 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=429  $PIN_XY=4118,444,4088,429,4058,444 $DEVICE_ID=1003
MM41 4 24 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=169  $PIN_XY=4118,154,4088,169,4058,154 $DEVICE_ID=1003
MM42 2 22 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=-495  $PIN_XY=4118,-480,4088,-495,4058,-480 $DEVICE_ID=1003
MM43 2 34 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=-755  $PIN_XY=4118,-770,4088,-755,4058,-770 $DEVICE_ID=1003
MM44 26 25 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=1353  $PIN_XY=3950,1368,3920,1353,3890,1368 $DEVICE_ID=1003
MM45 32 21 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=1093  $PIN_XY=3950,1078,3920,1093,3890,1078 $DEVICE_ID=1003
MM46 31 36 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=429  $PIN_XY=3950,444,3920,429,3890,444 $DEVICE_ID=1003
MM47 30 24 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=169  $PIN_XY=3950,154,3920,169,3890,154 $DEVICE_ID=1003
MM48 29 22 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=-495  $PIN_XY=3950,-480,3920,-495,3890,-480 $DEVICE_ID=1003
MM49 28 34 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=-755  $PIN_XY=3950,-770,3920,-755,3890,-770 $DEVICE_ID=1003
MM50 7 25 26 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=1454  $PIN_XY=3782,1368,3752,1454,3722,1368 $DEVICE_ID=1003
MM51 7 21 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=992  $PIN_XY=3782,1078,3752,992,3722,1078 $DEVICE_ID=1003
MM52 4 36 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=530  $PIN_XY=3782,444,3752,530,3722,444 $DEVICE_ID=1003
MM53 4 24 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=68  $PIN_XY=3782,154,3752,68,3722,154 $DEVICE_ID=1003
MM54 2 22 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=-394  $PIN_XY=3782,-480,3752,-394,3722,-480 $DEVICE_ID=1003
MM55 2 34 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=-856  $PIN_XY=3782,-770,3752,-856,3722,-770 $DEVICE_ID=1003
MM56 26 25 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=1454  $PIN_XY=3614,1368,3584,1454,3554,1368 $DEVICE_ID=1003
MM57 32 21 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=992  $PIN_XY=3614,1078,3584,992,3554,1078 $DEVICE_ID=1003
MM58 31 36 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=530  $PIN_XY=3614,444,3584,530,3554,444 $DEVICE_ID=1003
MM59 30 24 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=68  $PIN_XY=3614,154,3584,68,3554,154 $DEVICE_ID=1003
MM60 29 22 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-394  $PIN_XY=3614,-480,3584,-394,3554,-480 $DEVICE_ID=1003
MM61 28 34 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-856  $PIN_XY=3614,-770,3584,-856,3554,-770 $DEVICE_ID=1003
MM62 7 12 50 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=971  $PIN_XY=3278,1078,3248,971,3218,1078 $DEVICE_ID=1003
MM63 4 17 49 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=551  $PIN_XY=3278,444,3248,551,3218,444 $DEVICE_ID=1003
MM64 2 11 48 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=-877  $PIN_XY=3278,-770,3248,-877,3218,-770 $DEVICE_ID=1003
MM65 7 20 25 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=1454  $PIN_XY=3110,1368,3080,1454,3050,1368 $DEVICE_ID=1003
MM66 50 20 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=992  $PIN_XY=3110,1078,3080,992,3050,1078 $DEVICE_ID=1003
MM67 49 20 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=530  $PIN_XY=3110,444,3080,530,3050,444 $DEVICE_ID=1003
MM68 4 20 24 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=68  $PIN_XY=3110,154,3080,68,3050,154 $DEVICE_ID=1003
MM69 2 20 22 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=-394  $PIN_XY=3110,-480,3080,-394,3050,-480 $DEVICE_ID=1003
MM70 48 20 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=-856  $PIN_XY=3110,-770,3080,-856,3050,-770 $DEVICE_ID=1003
MM71 25 14 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=1475  $PIN_XY=2942,1368,2912,1475,2882,1368 $DEVICE_ID=1003
MM72 24 16 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=47  $PIN_XY=2942,154,2912,47,2882,154 $DEVICE_ID=1003
MM73 22 13 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=-373  $PIN_XY=2942,-480,2912,-373,2882,-480 $DEVICE_ID=1003
MM74 7 19 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2576 $Y=1072  $PIN_XY=2606,1078,2576,1072,2546,1078 $DEVICE_ID=1003
MM75 20 19 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2408 $Y=992  $PIN_XY=2438,1078,2408,992,2378,1078 $DEVICE_ID=1003
MM76 7 12 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2072 $Y=1454  $PIN_XY=2102,1368,2072,1454,2042,1368 $DEVICE_ID=1003
MM77 4 13 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2072 $Y=154  $PIN_XY=2102,154,2072,154,2042,154 $DEVICE_ID=1003
MM78 2 11 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2072 $Y=-394  $PIN_XY=2102,-480,2072,-394,2042,-480 $DEVICE_ID=1003
MM79 17 12 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1904 $Y=1374  $PIN_XY=1934,1368,1904,1374,1874,1368 $DEVICE_ID=1003
MM80 16 13 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1904 $Y=68  $PIN_XY=1934,154,1904,68,1874,154 $DEVICE_ID=1003
MM81 15 11 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1904 $Y=-474  $PIN_XY=1934,-480,1904,-474,1874,-480 $DEVICE_ID=1003
MM82 7 54 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1568 $Y=1374  $PIN_XY=1598,1368,1568,1374,1538,1368 $DEVICE_ID=1003
MM83 4 52 13 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1568 $Y=148  $PIN_XY=1598,154,1568,148,1538,154 $DEVICE_ID=1003
MM84 2 53 11 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1568 $Y=-474  $PIN_XY=1598,-480,1568,-474,1538,-480 $DEVICE_ID=1003
MM85 12 54 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1400 $Y=1475  $PIN_XY=1430,1368,1400,1475,1370,1368 $DEVICE_ID=1003
MM86 13 52 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1400 $Y=47  $PIN_XY=1430,154,1400,47,1370,154 $DEVICE_ID=1003
MM87 11 53 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1400 $Y=-373  $PIN_XY=1430,-480,1400,-373,1370,-480 $DEVICE_ID=1003
MM88 7 19 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=896 $Y=1475  $PIN_XY=926,1368,896,1475,866,1368 $DEVICE_ID=1003
MM89 4 51 52 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=896 $Y=47  $PIN_XY=926,154,896,47,866,154 $DEVICE_ID=1003
MM90 2 19 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=896 $Y=-373  $PIN_XY=926,-480,896,-373,866,-480 $DEVICE_ID=1003
MM91 54 38 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=728 $Y=1475  $PIN_XY=758,1368,728,1475,698,1368 $DEVICE_ID=1003
MM92 52 37 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=728 $Y=47  $PIN_XY=758,154,728,47,698,154 $DEVICE_ID=1003
MM93 53 37 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=728 $Y=-373  $PIN_XY=758,-480,728,-373,698,-480 $DEVICE_ID=1003
MM94 4 19 51 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=392 $Y=148  $PIN_XY=422,154,392,148,362,154 $DEVICE_ID=1003
MM95 51 19 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=224 $Y=68  $PIN_XY=254,154,224,68,194,154 $DEVICE_ID=1003
XX30BB92C5933 3 2 15 11 41 43 inv $T=2294 -100 0 180 $X=1682 $Y=-690
XX30BB92C5934 3 4 16 13 41 44 inv $T=1682 -226 0 0 $X=1682 $Y=-226
XX30BB92C5935 10 7 20 19 40 46 inv $T=2186 698 0 0 $X=2186 $Y=698
XX30BB92C5936 8 7 17 12 42 46 inv $T=2294 1748 0 180 $X=1682 $Y=1158
XX30BB92C5937 8 9 18 14 42 47 inv $T=1682 1622 0 0 $X=1682 $Y=1622
XX30BB92C5938 5 2 34 20 11 48 39 43 nor $T=4098 -1152 1 180 $X=2690 $Y=-1150
XX30BB92C5939 5 6 35 20 15 59 39 45 nor $T=4098 -1022 0 180 $X=2690 $Y=-1613
XX30BB92C5940 10 4 36 20 17 49 40 44 nor $T=4098 826 0 180 $X=2690 $Y=234
XX30BB92C5941 10 7 21 20 12 50 40 46 nor $T=4098 696 1 180 $X=2690 $Y=698
XX30BB92C5942 3 2 22 13 20 55 41 43 nand $T=2272 128 1 0 $X=2690 $Y=-690
XX30BB92C5943 3 4 24 16 20 56 41 44 nand $T=2272 -454 0 0 $X=2690 $Y=-226
XX30BB92C5944 8 7 25 14 20 57 42 46 nand $T=2272 1976 1 0 $X=2690 $Y=1158
XX30BB92C5945 8 9 23 18 20 58 42 47 nand $T=2272 1394 0 0 $X=2690 $Y=1622
XX30BB92C5946 3 2 4 19 51 37 53 52 11 13 41 
+	43 44 Demux $T=2 -688 0 0 $X=2 $Y=-690
XX30BB92C5947 8 7 9 19 60 38 54 61 12 14 42 
+	46 47 Demux $T=2 1160 0 0 $X=2 $Y=1158
XX30BB92C5948 3 4 30 24 41 44 invx4 $T=3338 -226 0 0 $X=3362 $Y=-226
XX30BB92C5949 10 4 31 36 40 44 invx4 $T=3338 824 1 0 $X=3362 $Y=234
XX30BB92C5950 5 6 27 35 39 45 invx4 $T=3338 -1024 1 0 $X=3362 $Y=-1613
XX30BB92C5951 3 2 29 22 41 43 invx4 $T=3338 -100 1 0 $X=3362 $Y=-690
XX30BB92C5952 5 2 28 34 39 43 invx4 $T=3338 -1150 0 0 $X=3362 $Y=-1150
XX30BB92C5953 8 9 33 23 42 47 invx4 $T=3338 1622 0 0 $X=3362 $Y=1622
XX30BB92C5954 8 7 26 25 42 46 invx4 $T=3338 1748 1 0 $X=3362 $Y=1158
XX30BB92C5955 10 7 32 21 40 46 invx4 $T=3338 698 0 0 $X=3362 $Y=698
XX30BB92C5956 5 6 _GENERATED_63 _GENERATED_62 39 45 sram_filler $T=-2 -1024 1 0 $X=2 $Y=-1613
XX30BB92C5957 5 6 _GENERATED_64 5 39 45 sram_filler $T=334 -1024 1 0 $X=338 $Y=-1613
XX30BB92C5958 5 6 6 _GENERATED_65 39 45 sram_filler $T=502 -1024 1 0 $X=506 $Y=-1613
XX30BB92C5959 5 2 _GENERATED_66 5 39 43 sram_filler $T=-2 -1150 0 0 $X=2 $Y=-1150
XX30BB92C5960 5 2 2 _GENERATED_67 39 43 sram_filler $T=166 -1150 0 0 $X=170 $Y=-1150
XX30BB92C5961 5 2 _GENERATED_69 _GENERATED_68 39 43 sram_filler $T=502 -1150 0 0 $X=506 $Y=-1150
XX30BB92C5962 5 6 6 _GENERATED_70 39 45 sram_filler $T=1342 -1024 1 0 $X=1346 $Y=-1613
XX30BB92C5963 5 6 _GENERATED_71 5 39 45 sram_filler $T=1174 -1024 1 0 $X=1178 $Y=-1613
XX30BB92C5964 5 6 _GENERATED_73 _GENERATED_72 39 45 sram_filler $T=838 -1024 1 0 $X=842 $Y=-1613
XX30BB92C5965 5 2 2 _GENERATED_74 39 43 sram_filler $T=1342 -1150 0 0 $X=1346 $Y=-1150
XX30BB92C5966 5 2 _GENERATED_75 5 39 43 sram_filler $T=1174 -1150 0 0 $X=1178 $Y=-1150
XX30BB92C5967 5 2 _GENERATED_77 _GENERATED_76 39 43 sram_filler $T=838 -1150 0 0 $X=842 $Y=-1150
XX30BB92C5968 5 2 _GENERATED_79 _GENERATED_78 39 43 sram_filler $T=1678 -1150 0 0 $X=1682 $Y=-1150
XX30BB92C5969 5 6 _GENERATED_81 _GENERATED_80 39 45 sram_filler $T=2130 -1024 0 180 $X=1682 $Y=-1613
XX30BB92C5970 10 7 7 _GENERATED_82 40 46 sram_filler $T=1846 698 0 0 $X=1850 $Y=698
XX30BB92C5971 10 4 _GENERATED_83 10 40 44 sram_filler $T=2298 824 0 180 $X=1850 $Y=234
XX30BB92C5972 5 2 _GENERATED_85 _GENERATED_84 39 43 sram_filler $T=2014 -1150 0 0 $X=2018 $Y=-1150
XX30BB92C5973 5 6 _GENERATED_87 _GENERATED_86 39 45 sram_filler $T=2466 -1024 0 180 $X=2018 $Y=-1613
XX30BB92C5974 5 6 _GENERATED_89 _GENERATED_88 39 45 sram_filler $T=2802 -1024 0 180 $X=2354 $Y=-1613
XX30BB92C5975 5 2 _GENERATED_91 _GENERATED_90 39 43 sram_filler $T=2350 -1150 0 0 $X=2354 $Y=-1150
XX30BB92C5976 10 4 _GENERATED_93 _GENERATED_92 40 44 sram_filler $T=1794 824 0 180 $X=1346 $Y=234
XX30BB92C5977 10 4 _GENERATED_95 _GENERATED_94 40 44 sram_filler $T=1458 824 0 180 $X=1010 $Y=234
XX30BB92C5978 10 4 _GENERATED_97 _GENERATED_96 40 44 sram_filler $T=1122 824 0 180 $X=674 $Y=234
XX30BB92C5979 10 4 _GENERATED_99 _GENERATED_98 40 44 sram_filler $T=786 824 0 180 $X=338 $Y=234
XX30BB92C5980 10 4 _GENERATED_101 _GENERATED_100 40 44 sram_filler $T=450 824 0 180 $X=2 $Y=234
XX30BB92C5981 10 7 7 _GENERATED_102 40 46 sram_filler $T=1342 698 0 0 $X=1346 $Y=698
XX30BB92C5982 10 7 _GENERATED_103 10 40 46 sram_filler $T=1174 698 0 0 $X=1178 $Y=698
XX30BB92C5983 10 7 _GENERATED_105 _GENERATED_104 40 46 sram_filler $T=838 698 0 0 $X=842 $Y=698
XX30BB92C5984 10 7 7 _GENERATED_106 40 46 sram_filler $T=502 698 0 0 $X=506 $Y=698
XX30BB92C5985 10 7 _GENERATED_107 10 40 46 sram_filler $T=334 698 0 0 $X=338 $Y=698
XX30BB92C5986 10 7 _GENERATED_109 _GENERATED_108 40 46 sram_filler $T=-2 698 0 0 $X=2 $Y=698
XX30BB92C5987 3 2 _GENERATED_110 3 41 43 sram_filler $T=2802 -100 0 180 $X=2354 $Y=-690
XX30BB92C5988 3 2 2 _GENERATED_111 41 43 sram_filler $T=2634 -100 0 180 $X=2186 $Y=-690
XX30BB92C5989 3 4 _GENERATED_112 3 41 44 sram_filler $T=2182 -226 0 0 $X=2186 $Y=-226
XX30BB92C5990 3 4 4 _GENERATED_113 41 44 sram_filler $T=2350 -226 0 0 $X=2354 $Y=-226
XX30BB92C5991 10 4 _GENERATED_114 10 40 44 sram_filler $T=2802 824 0 180 $X=2354 $Y=234
XX30BB92C5992 10 4 4 _GENERATED_115 40 44 sram_filler $T=2634 824 0 180 $X=2186 $Y=234
XX30BB92C5993 8 7 _GENERATED_116 8 42 46 sram_filler $T=2802 1748 0 180 $X=2354 $Y=1158
XX30BB92C5994 8 7 7 _GENERATED_117 42 46 sram_filler $T=2634 1748 0 180 $X=2186 $Y=1158
XX30BB92C5995 8 9 9 _GENERATED_118 42 47 sram_filler $T=2350 1622 0 0 $X=2354 $Y=1622
XX30BB92C5996 8 9 _GENERATED_119 8 42 47 sram_filler $T=2182 1622 0 0 $X=2186 $Y=1622
XX30BB92C5997 10 7 _GENERATED_120 10 40 46 sram_filler $T=1678 698 0 0 $X=1682 $Y=698
XX30BB92C5998 10 4 4 _GENERATED_121 40 44 sram_filler $T=2130 824 0 180 $X=1682 $Y=234
.ends agen_unit
.subckt Write_Driver 2 3 4 6 7 8 9 10 11 12 13
+	14 15 16 17 18 19 20 21 22 23 24
+	25
MM1 3 25 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2386 $Y=852  $PIN_XY=2416,936,2386,852,2356,936 $DEVICE_ID=1001
MM2 10 25 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2218 $Y=852  $PIN_XY=2248,936,2218,852,2188,936 $DEVICE_ID=1001
MM3 3 8 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1546 $Y=1293  $PIN_XY=1576,1230,1546,1293,1516,1230 $DEVICE_ID=1001
MM4 3 7 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1546 $Y=873  $PIN_XY=1576,936,1546,873,1516,936 $DEVICE_ID=1001
MM5 9 8 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1378 $Y=1293  $PIN_XY=1408,1230,1378,1293,1348,1230 $DEVICE_ID=1001
MM6 25 7 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1378 $Y=852  $PIN_XY=1408,936,1378,852,1348,936 $DEVICE_ID=1001
MM7 8 12 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=874 $Y=1293  $PIN_XY=904,1230,874,1293,844,1230 $DEVICE_ID=1001
MM8 7 11 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=874 $Y=852  $PIN_XY=904,936,874,852,844,936 $DEVICE_ID=1001
MM9 12 6 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=370 $Y=1293  $PIN_XY=400,1230,370,1293,340,1230 $DEVICE_ID=1001
MM10 11 6 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=370 $Y=852  $PIN_XY=400,936,370,852,340,936 $DEVICE_ID=1001
XX30BB92C51031 2 3 10 25 7 21 22 23 buffer_highdrive $T=1154 1144 1 0 $X=1156 $Y=556
XX30BB92C51032 3 2 11 7 6 22 23 buffer $T=68 1148 1 0 $X=148 $Y=556
XX30BB92C51033 3 4 12 8 6 22 24 buffer $T=68 1018 0 0 $X=148 $Y=1020
XX30BB92C51034 3 2 17 18 22 23 sram_filler $T=3284 1146 0 180 $X=2836 $Y=556
XX30BB92C51035 3 4 19 20 22 24 sram_filler $T=3284 1020 1 180 $X=2836 $Y=1020
XX30BB92C51036 3 4 _GENERATED_26 5 22 24 sram_filler $T=2948 1020 1 180 $X=2500 $Y=1020
XX30BB92C51037 3 4 _GENERATED_27 5 22 24 sram_filler $T=2328 1020 0 0 $X=2332 $Y=1020
XX30BB92C51038 3 4 _GENERATED_29 _GENERATED_28 22 24 sram_filler $T=1992 1020 0 0 $X=1996 $Y=1020
XX30BB92C51039 3 4 9 8 22 24 invx4 $T=1132 1020 0 0 $X=1156 $Y=1020
.ends Write_Driver

* Hierarchy Level 0

* Top of hierarchy  cell=integration
.subckt integration GND! VDD! Q<1> Q<0> Q<2> Q<3> 8 9 10 11 12
+	13 14 15 16 17 18 19 20 21 22 23
+	24 25 26 27 WS1 WS1BAR 63 64 65 66 67
+	68 69 70 71 72 73 74 75 76 77 78
+	79 80 WS0 82 83 WENB 85 86 87 WS0BAR 89
+	90 91 92 93 94 CLK 96 97 98 99 100
+	A<4> A<3> 103 104 105 106 107 108 D<0> D<1> D<2>
+	D<3> 113 A<1> A<0> A<2>
MM1 GND! 454 256 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=14616  $PIN_XY=18174,14700,18144,14616,18114,14700 $DEVICE_ID=1001
MM2 27 108 454 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=14067  $PIN_XY=18174,14070,18144,14067,18114,14070 $DEVICE_ID=1001
MM3 GND! 452 251 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=13692  $PIN_XY=18174,13776,18144,13692,18114,13776 $DEVICE_ID=1001
MM4 27 107 452 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=13143  $PIN_XY=18174,13146,18144,13143,18114,13146 $DEVICE_ID=1001
MM5 GND! 447 245 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=12768  $PIN_XY=18174,12852,18144,12768,18114,12852 $DEVICE_ID=1001
MM6 27 106 447 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=12219  $PIN_XY=18174,12222,18144,12219,18114,12222 $DEVICE_ID=1001
MM7 GND! 405 242 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=11844  $PIN_XY=18174,11928,18144,11844,18114,11928 $DEVICE_ID=1001
MM8 256 108 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=14703  $PIN_XY=18006,14700,17976,14703,17946,14700 $DEVICE_ID=1001
MM9 454 256 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=14154  $PIN_XY=18006,14070,17976,14154,17946,14070 $DEVICE_ID=1001
MM10 251 107 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=13779  $PIN_XY=18006,13776,17976,13779,17946,13776 $DEVICE_ID=1001
MM11 452 251 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=13230  $PIN_XY=18006,13146,17976,13230,17946,13146 $DEVICE_ID=1001
MM12 245 106 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=12855  $PIN_XY=18006,12852,17976,12855,17946,12852 $DEVICE_ID=1001
MM13 447 245 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=12306  $PIN_XY=18006,12222,17976,12306,17946,12222 $DEVICE_ID=1001
MM14 242 105 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=11931  $PIN_XY=18006,11928,17976,11931,17946,11928 $DEVICE_ID=1001
MM15 GND! 455 255 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=14616  $PIN_XY=17502,14700,17472,14616,17442,14700 $DEVICE_ID=1001
MM16 26 108 455 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=14067  $PIN_XY=17502,14070,17472,14067,17442,14070 $DEVICE_ID=1001
MM17 GND! 451 250 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=13692  $PIN_XY=17502,13776,17472,13692,17442,13776 $DEVICE_ID=1001
MM18 26 107 451 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=13143  $PIN_XY=17502,13146,17472,13143,17442,13146 $DEVICE_ID=1001
MM19 GND! 446 246 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=12768  $PIN_XY=17502,12852,17472,12768,17442,12852 $DEVICE_ID=1001
MM20 26 106 446 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=12219  $PIN_XY=17502,12222,17472,12219,17442,12222 $DEVICE_ID=1001
MM21 GND! 406 243 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=11844  $PIN_XY=17502,11928,17472,11844,17442,11928 $DEVICE_ID=1001
MM22 255 108 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=14703  $PIN_XY=17334,14700,17304,14703,17274,14700 $DEVICE_ID=1001
MM23 455 255 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=14154  $PIN_XY=17334,14070,17304,14154,17274,14070 $DEVICE_ID=1001
MM24 250 107 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=13779  $PIN_XY=17334,13776,17304,13779,17274,13776 $DEVICE_ID=1001
MM25 451 250 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=13230  $PIN_XY=17334,13146,17304,13230,17274,13146 $DEVICE_ID=1001
MM26 246 106 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=12855  $PIN_XY=17334,12852,17304,12855,17274,12852 $DEVICE_ID=1001
MM27 446 246 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=12306  $PIN_XY=17334,12222,17304,12306,17274,12222 $DEVICE_ID=1001
MM28 243 105 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=11931  $PIN_XY=17334,11928,17304,11931,17274,11928 $DEVICE_ID=1001
MM29 GND! 456 254 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=14616  $PIN_XY=16830,14700,16800,14616,16770,14700 $DEVICE_ID=1001
MM30 25 108 456 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=14067  $PIN_XY=16830,14070,16800,14067,16770,14070 $DEVICE_ID=1001
MM31 GND! 450 249 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=13692  $PIN_XY=16830,13776,16800,13692,16770,13776 $DEVICE_ID=1001
MM32 25 107 450 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=13143  $PIN_XY=16830,13146,16800,13143,16770,13146 $DEVICE_ID=1001
MM33 GND! 445 247 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=12768  $PIN_XY=16830,12852,16800,12768,16770,12852 $DEVICE_ID=1001
MM34 25 106 445 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=12219  $PIN_XY=16830,12222,16800,12219,16770,12222 $DEVICE_ID=1001
MM35 GND! 407 244 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=11844  $PIN_XY=16830,11928,16800,11844,16770,11928 $DEVICE_ID=1001
MM36 254 108 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=14703  $PIN_XY=16662,14700,16632,14703,16602,14700 $DEVICE_ID=1001
MM37 456 254 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=14154  $PIN_XY=16662,14070,16632,14154,16602,14070 $DEVICE_ID=1001
MM38 249 107 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=13779  $PIN_XY=16662,13776,16632,13779,16602,13776 $DEVICE_ID=1001
MM39 450 249 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=13230  $PIN_XY=16662,13146,16632,13230,16602,13146 $DEVICE_ID=1001
MM40 247 106 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=12855  $PIN_XY=16662,12852,16632,12855,16602,12852 $DEVICE_ID=1001
MM41 445 247 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=12306  $PIN_XY=16662,12222,16632,12306,16602,12222 $DEVICE_ID=1001
MM42 244 105 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=11931  $PIN_XY=16662,11928,16632,11931,16602,11928 $DEVICE_ID=1001
MM43 27 105 405 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=11295  $PIN_XY=18174,11298,18144,11295,18114,11298 $DEVICE_ID=1001
MM44 GND! 402 240 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=10920  $PIN_XY=18174,11004,18144,10920,18114,11004 $DEVICE_ID=1001
MM45 27 104 402 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=10371  $PIN_XY=18174,10374,18144,10371,18114,10374 $DEVICE_ID=1001
MM46 GND! 400 170 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=9996  $PIN_XY=18174,10080,18144,9996,18114,10080 $DEVICE_ID=1001
MM47 27 103 400 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=9447  $PIN_XY=18174,9450,18144,9447,18114,9450 $DEVICE_ID=1001
MM48 GND! 357 169 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=9072  $PIN_XY=18174,9156,18144,9072,18114,9156 $DEVICE_ID=1001
MM49 27 99 357 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=8523  $PIN_XY=18174,8526,18144,8523,18114,8526 $DEVICE_ID=1001
MM50 405 242 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=11382  $PIN_XY=18006,11298,17976,11382,17946,11298 $DEVICE_ID=1001
MM51 240 104 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=11007  $PIN_XY=18006,11004,17976,11007,17946,11004 $DEVICE_ID=1001
MM52 402 240 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=10458  $PIN_XY=18006,10374,17976,10458,17946,10374 $DEVICE_ID=1001
MM53 170 103 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=10083  $PIN_XY=18006,10080,17976,10083,17946,10080 $DEVICE_ID=1001
MM54 400 170 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=9534  $PIN_XY=18006,9450,17976,9534,17946,9450 $DEVICE_ID=1001
MM55 169 99 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=9159  $PIN_XY=18006,9156,17976,9159,17946,9156 $DEVICE_ID=1001
MM56 357 169 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=8610  $PIN_XY=18006,8526,17976,8610,17946,8526 $DEVICE_ID=1001
MM57 26 105 406 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=11295  $PIN_XY=17502,11298,17472,11295,17442,11298 $DEVICE_ID=1001
MM58 GND! 403 239 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=10920  $PIN_XY=17502,11004,17472,10920,17442,11004 $DEVICE_ID=1001
MM59 26 104 403 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=10371  $PIN_XY=17502,10374,17472,10371,17442,10374 $DEVICE_ID=1001
MM60 GND! 399 172 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=9996  $PIN_XY=17502,10080,17472,9996,17442,10080 $DEVICE_ID=1001
MM61 26 103 399 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=9447  $PIN_XY=17502,9450,17472,9447,17442,9450 $DEVICE_ID=1001
MM62 GND! 358 171 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=9072  $PIN_XY=17502,9156,17472,9072,17442,9156 $DEVICE_ID=1001
MM63 26 99 358 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=8523  $PIN_XY=17502,8526,17472,8523,17442,8526 $DEVICE_ID=1001
MM64 406 243 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=11382  $PIN_XY=17334,11298,17304,11382,17274,11298 $DEVICE_ID=1001
MM65 239 104 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=11007  $PIN_XY=17334,11004,17304,11007,17274,11004 $DEVICE_ID=1001
MM66 403 239 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=10458  $PIN_XY=17334,10374,17304,10458,17274,10374 $DEVICE_ID=1001
MM67 172 103 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=10083  $PIN_XY=17334,10080,17304,10083,17274,10080 $DEVICE_ID=1001
MM68 399 172 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=9534  $PIN_XY=17334,9450,17304,9534,17274,9450 $DEVICE_ID=1001
MM69 171 99 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=9159  $PIN_XY=17334,9156,17304,9159,17274,9156 $DEVICE_ID=1001
MM70 358 171 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=8610  $PIN_XY=17334,8526,17304,8610,17274,8526 $DEVICE_ID=1001
MM71 25 105 407 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=11295  $PIN_XY=16830,11298,16800,11295,16770,11298 $DEVICE_ID=1001
MM72 GND! 404 238 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=10920  $PIN_XY=16830,11004,16800,10920,16770,11004 $DEVICE_ID=1001
MM73 25 104 404 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=10371  $PIN_XY=16830,10374,16800,10371,16770,10374 $DEVICE_ID=1001
MM74 GND! 398 174 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=9996  $PIN_XY=16830,10080,16800,9996,16770,10080 $DEVICE_ID=1001
MM75 25 103 398 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=9447  $PIN_XY=16830,9450,16800,9447,16770,9450 $DEVICE_ID=1001
MM76 GND! 359 173 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=9072  $PIN_XY=16830,9156,16800,9072,16770,9156 $DEVICE_ID=1001
MM77 25 99 359 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=8523  $PIN_XY=16830,8526,16800,8523,16770,8526 $DEVICE_ID=1001
MM78 407 244 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=11382  $PIN_XY=16662,11298,16632,11382,16602,11298 $DEVICE_ID=1001
MM79 238 104 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=11007  $PIN_XY=16662,11004,16632,11007,16602,11004 $DEVICE_ID=1001
MM80 404 238 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=10458  $PIN_XY=16662,10374,16632,10458,16602,10374 $DEVICE_ID=1001
MM81 174 103 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=10083  $PIN_XY=16662,10080,16632,10083,16602,10080 $DEVICE_ID=1001
MM82 398 174 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=9534  $PIN_XY=16662,9450,16632,9534,16602,9450 $DEVICE_ID=1001
MM83 173 99 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=9159  $PIN_XY=16662,9156,16632,9159,16602,9156 $DEVICE_ID=1001
MM84 359 173 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=8610  $PIN_XY=16662,8526,16632,8610,16602,8526 $DEVICE_ID=1001
MM85 GND! 453 253 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=14616  $PIN_XY=16158,14700,16128,14616,16098,14700 $DEVICE_ID=1001
MM86 23 108 453 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=14067  $PIN_XY=16158,14070,16128,14067,16098,14070 $DEVICE_ID=1001
MM87 GND! 449 252 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=13692  $PIN_XY=16158,13776,16128,13692,16098,13776 $DEVICE_ID=1001
MM88 23 107 449 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=13143  $PIN_XY=16158,13146,16128,13143,16098,13146 $DEVICE_ID=1001
MM89 GND! 448 248 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=12768  $PIN_XY=16158,12852,16128,12768,16098,12852 $DEVICE_ID=1001
MM90 23 106 448 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=12219  $PIN_XY=16158,12222,16128,12219,16098,12222 $DEVICE_ID=1001
MM91 GND! 408 241 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=11844  $PIN_XY=16158,11928,16128,11844,16098,11928 $DEVICE_ID=1001
MM92 253 108 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=14703  $PIN_XY=15990,14700,15960,14703,15930,14700 $DEVICE_ID=1001
MM93 453 253 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=14154  $PIN_XY=15990,14070,15960,14154,15930,14070 $DEVICE_ID=1001
MM94 252 107 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=13779  $PIN_XY=15990,13776,15960,13779,15930,13776 $DEVICE_ID=1001
MM95 449 252 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=13230  $PIN_XY=15990,13146,15960,13230,15930,13146 $DEVICE_ID=1001
MM96 248 106 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=12855  $PIN_XY=15990,12852,15960,12855,15930,12852 $DEVICE_ID=1001
MM97 448 248 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=12306  $PIN_XY=15990,12222,15960,12306,15930,12222 $DEVICE_ID=1001
MM98 241 105 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=11931  $PIN_XY=15990,11928,15960,11931,15930,11928 $DEVICE_ID=1001
MM99 GND! 457 217 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=14616  $PIN_XY=15150,14700,15120,14616,15090,14700 $DEVICE_ID=1001
MM100 22 108 457 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=14067  $PIN_XY=15150,14070,15120,14067,15090,14070 $DEVICE_ID=1001
MM101 GND! 458 218 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=13692  $PIN_XY=15150,13776,15120,13692,15090,13776 $DEVICE_ID=1001
MM102 22 107 458 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=13143  $PIN_XY=15150,13146,15120,13143,15090,13146 $DEVICE_ID=1001
MM103 GND! 459 219 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=12768  $PIN_XY=15150,12852,15120,12768,15090,12852 $DEVICE_ID=1001
MM104 22 106 459 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=12219  $PIN_XY=15150,12222,15120,12219,15090,12222 $DEVICE_ID=1001
MM105 GND! 409 220 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=11844  $PIN_XY=15150,11928,15120,11844,15090,11928 $DEVICE_ID=1001
MM106 217 108 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=14703  $PIN_XY=14982,14700,14952,14703,14922,14700 $DEVICE_ID=1001
MM107 457 217 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=14154  $PIN_XY=14982,14070,14952,14154,14922,14070 $DEVICE_ID=1001
MM108 218 107 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=13779  $PIN_XY=14982,13776,14952,13779,14922,13776 $DEVICE_ID=1001
MM109 458 218 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=13230  $PIN_XY=14982,13146,14952,13230,14922,13146 $DEVICE_ID=1001
MM110 219 106 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=12855  $PIN_XY=14982,12852,14952,12855,14922,12852 $DEVICE_ID=1001
MM111 459 219 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=12306  $PIN_XY=14982,12222,14952,12306,14922,12222 $DEVICE_ID=1001
MM112 220 105 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=11931  $PIN_XY=14982,11928,14952,11931,14922,11928 $DEVICE_ID=1001
MM113 GND! 461 223 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=14616  $PIN_XY=14478,14700,14448,14616,14418,14700 $DEVICE_ID=1001
MM114 18 108 461 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=14067  $PIN_XY=14478,14070,14448,14067,14418,14070 $DEVICE_ID=1001
MM115 GND! 463 225 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=13692  $PIN_XY=14478,13776,14448,13692,14418,13776 $DEVICE_ID=1001
MM116 18 107 463 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=13143  $PIN_XY=14478,13146,14448,13143,14418,13146 $DEVICE_ID=1001
MM117 GND! 467 229 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=12768  $PIN_XY=14478,12852,14448,12768,14418,12852 $DEVICE_ID=1001
MM118 18 106 467 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=12219  $PIN_XY=14478,12222,14448,12219,14418,12222 $DEVICE_ID=1001
MM119 GND! 414 233 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=11844  $PIN_XY=14478,11928,14448,11844,14418,11928 $DEVICE_ID=1001
MM120 223 108 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=14703  $PIN_XY=14310,14700,14280,14703,14250,14700 $DEVICE_ID=1001
MM121 461 223 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=14154  $PIN_XY=14310,14070,14280,14154,14250,14070 $DEVICE_ID=1001
MM122 225 107 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=13779  $PIN_XY=14310,13776,14280,13779,14250,13776 $DEVICE_ID=1001
MM123 463 225 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=13230  $PIN_XY=14310,13146,14280,13230,14250,13146 $DEVICE_ID=1001
MM124 229 106 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=12855  $PIN_XY=14310,12852,14280,12855,14250,12852 $DEVICE_ID=1001
MM125 467 229 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=12306  $PIN_XY=14310,12222,14280,12306,14250,12222 $DEVICE_ID=1001
MM126 233 105 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=11931  $PIN_XY=14310,11928,14280,11931,14250,11928 $DEVICE_ID=1001
MM127 23 105 408 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=11295  $PIN_XY=16158,11298,16128,11295,16098,11298 $DEVICE_ID=1001
MM128 GND! 401 237 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=10920  $PIN_XY=16158,11004,16128,10920,16098,11004 $DEVICE_ID=1001
MM129 23 104 401 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=10371  $PIN_XY=16158,10374,16128,10371,16098,10374 $DEVICE_ID=1001
MM130 GND! 397 176 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=9996  $PIN_XY=16158,10080,16128,9996,16098,10080 $DEVICE_ID=1001
MM131 23 103 397 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=9447  $PIN_XY=16158,9450,16128,9447,16098,9450 $DEVICE_ID=1001
MM132 GND! 360 175 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=9072  $PIN_XY=16158,9156,16128,9072,16098,9156 $DEVICE_ID=1001
MM133 23 99 360 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=8523  $PIN_XY=16158,8526,16128,8523,16098,8526 $DEVICE_ID=1001
MM134 408 241 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=11382  $PIN_XY=15990,11298,15960,11382,15930,11298 $DEVICE_ID=1001
MM135 237 104 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=11007  $PIN_XY=15990,11004,15960,11007,15930,11004 $DEVICE_ID=1001
MM136 401 237 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=10458  $PIN_XY=15990,10374,15960,10458,15930,10374 $DEVICE_ID=1001
MM137 176 103 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=10083  $PIN_XY=15990,10080,15960,10083,15930,10080 $DEVICE_ID=1001
MM138 397 176 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=9534  $PIN_XY=15990,9450,15960,9534,15930,9450 $DEVICE_ID=1001
MM139 175 99 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=9159  $PIN_XY=15990,9156,15960,9159,15930,9156 $DEVICE_ID=1001
MM140 360 175 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=8610  $PIN_XY=15990,8526,15960,8610,15930,8526 $DEVICE_ID=1001
MM141 22 105 409 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=11295  $PIN_XY=15150,11298,15120,11295,15090,11298 $DEVICE_ID=1001
MM142 GND! 410 221 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=10920  $PIN_XY=15150,11004,15120,10920,15090,11004 $DEVICE_ID=1001
MM143 22 104 410 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=10371  $PIN_XY=15150,10374,15120,10371,15090,10374 $DEVICE_ID=1001
MM144 GND! 411 158 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=9996  $PIN_XY=15150,10080,15120,9996,15090,10080 $DEVICE_ID=1001
MM145 22 103 411 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=9447  $PIN_XY=15150,9450,15120,9447,15090,9450 $DEVICE_ID=1001
MM146 GND! 361 157 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=9072  $PIN_XY=15150,9156,15120,9072,15090,9156 $DEVICE_ID=1001
MM147 22 99 361 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=8523  $PIN_XY=15150,8526,15120,8523,15090,8526 $DEVICE_ID=1001
MM148 409 220 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=11382  $PIN_XY=14982,11298,14952,11382,14922,11298 $DEVICE_ID=1001
MM149 221 104 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=11007  $PIN_XY=14982,11004,14952,11007,14922,11004 $DEVICE_ID=1001
MM150 410 221 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=10458  $PIN_XY=14982,10374,14952,10458,14922,10374 $DEVICE_ID=1001
MM151 158 103 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=10083  $PIN_XY=14982,10080,14952,10083,14922,10080 $DEVICE_ID=1001
MM152 411 158 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=9534  $PIN_XY=14982,9450,14952,9534,14922,9450 $DEVICE_ID=1001
MM153 157 99 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=9159  $PIN_XY=14982,9156,14952,9159,14922,9156 $DEVICE_ID=1001
MM154 361 157 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=8610  $PIN_XY=14982,8526,14952,8610,14922,8526 $DEVICE_ID=1001
MM155 18 105 414 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=11295  $PIN_XY=14478,11298,14448,11295,14418,11298 $DEVICE_ID=1001
MM156 GND! 416 235 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=10920  $PIN_XY=14478,11004,14448,10920,14418,11004 $DEVICE_ID=1001
MM157 18 104 416 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=10371  $PIN_XY=14478,10374,14448,10371,14418,10374 $DEVICE_ID=1001
MM158 GND! 418 164 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=9996  $PIN_XY=14478,10080,14448,9996,14418,10080 $DEVICE_ID=1001
MM159 18 103 418 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=9447  $PIN_XY=14478,9450,14448,9447,14418,9450 $DEVICE_ID=1001
MM160 GND! 368 163 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=9072  $PIN_XY=14478,9156,14448,9072,14418,9156 $DEVICE_ID=1001
MM161 18 99 368 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=8523  $PIN_XY=14478,8526,14448,8523,14418,8526 $DEVICE_ID=1001
MM162 414 233 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=11382  $PIN_XY=14310,11298,14280,11382,14250,11298 $DEVICE_ID=1001
MM163 235 104 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=11007  $PIN_XY=14310,11004,14280,11007,14250,11004 $DEVICE_ID=1001
MM164 416 235 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=10458  $PIN_XY=14310,10374,14280,10458,14250,10374 $DEVICE_ID=1001
MM165 164 103 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=10083  $PIN_XY=14310,10080,14280,10083,14250,10080 $DEVICE_ID=1001
MM166 418 164 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=9534  $PIN_XY=14310,9450,14280,9534,14250,9450 $DEVICE_ID=1001
MM167 163 99 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=9159  $PIN_XY=14310,9156,14280,9159,14250,9156 $DEVICE_ID=1001
MM168 368 163 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=8610  $PIN_XY=14310,8526,14280,8610,14250,8526 $DEVICE_ID=1001
MM169 GND! 460 222 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=14616  $PIN_XY=13806,14700,13776,14616,13746,14700 $DEVICE_ID=1001
MM170 20 108 460 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=14067  $PIN_XY=13806,14070,13776,14067,13746,14070 $DEVICE_ID=1001
MM171 GND! 464 226 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=13692  $PIN_XY=13806,13776,13776,13692,13746,13776 $DEVICE_ID=1001
MM172 20 107 464 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=13143  $PIN_XY=13806,13146,13776,13143,13746,13146 $DEVICE_ID=1001
MM173 GND! 468 230 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=12768  $PIN_XY=13806,12852,13776,12768,13746,12852 $DEVICE_ID=1001
MM174 20 106 468 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=12219  $PIN_XY=13806,12222,13776,12219,13746,12222 $DEVICE_ID=1001
MM175 GND! 413 232 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=11844  $PIN_XY=13806,11928,13776,11844,13746,11928 $DEVICE_ID=1001
MM176 20 105 413 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=11295  $PIN_XY=13806,11298,13776,11295,13746,11298 $DEVICE_ID=1001
MM177 GND! 415 234 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=10920  $PIN_XY=13806,11004,13776,10920,13746,11004 $DEVICE_ID=1001
MM178 20 104 415 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=10371  $PIN_XY=13806,10374,13776,10371,13746,10374 $DEVICE_ID=1001
MM179 GND! 419 162 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=9996  $PIN_XY=13806,10080,13776,9996,13746,10080 $DEVICE_ID=1001
MM180 20 103 419 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=9447  $PIN_XY=13806,9450,13776,9447,13746,9450 $DEVICE_ID=1001
MM181 GND! 367 161 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=9072  $PIN_XY=13806,9156,13776,9072,13746,9156 $DEVICE_ID=1001
MM182 20 99 367 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=8523  $PIN_XY=13806,8526,13776,8523,13746,8526 $DEVICE_ID=1001
MM183 222 108 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=14703  $PIN_XY=13638,14700,13608,14703,13578,14700 $DEVICE_ID=1001
MM184 460 222 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=14154  $PIN_XY=13638,14070,13608,14154,13578,14070 $DEVICE_ID=1001
MM185 226 107 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=13779  $PIN_XY=13638,13776,13608,13779,13578,13776 $DEVICE_ID=1001
MM186 464 226 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=13230  $PIN_XY=13638,13146,13608,13230,13578,13146 $DEVICE_ID=1001
MM187 230 106 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=12855  $PIN_XY=13638,12852,13608,12855,13578,12852 $DEVICE_ID=1001
MM188 468 230 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=12306  $PIN_XY=13638,12222,13608,12306,13578,12222 $DEVICE_ID=1001
MM189 232 105 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=11931  $PIN_XY=13638,11928,13608,11931,13578,11928 $DEVICE_ID=1001
MM190 413 232 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=11382  $PIN_XY=13638,11298,13608,11382,13578,11298 $DEVICE_ID=1001
MM191 234 104 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=11007  $PIN_XY=13638,11004,13608,11007,13578,11004 $DEVICE_ID=1001
MM192 415 234 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=10458  $PIN_XY=13638,10374,13608,10458,13578,10374 $DEVICE_ID=1001
MM193 162 103 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=10083  $PIN_XY=13638,10080,13608,10083,13578,10080 $DEVICE_ID=1001
MM194 419 162 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=9534  $PIN_XY=13638,9450,13608,9534,13578,9450 $DEVICE_ID=1001
MM195 161 99 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=9159  $PIN_XY=13638,9156,13608,9159,13578,9156 $DEVICE_ID=1001
MM196 367 161 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=8610  $PIN_XY=13638,8526,13608,8610,13578,8526 $DEVICE_ID=1001
MM197 GND! 462 224 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=14616  $PIN_XY=13134,14700,13104,14616,13074,14700 $DEVICE_ID=1001
MM198 21 108 462 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=14067  $PIN_XY=13134,14070,13104,14067,13074,14070 $DEVICE_ID=1001
MM199 GND! 465 227 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=13692  $PIN_XY=13134,13776,13104,13692,13074,13776 $DEVICE_ID=1001
MM200 21 107 465 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=13143  $PIN_XY=13134,13146,13104,13143,13074,13146 $DEVICE_ID=1001
MM201 GND! 466 228 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=12768  $PIN_XY=13134,12852,13104,12768,13074,12852 $DEVICE_ID=1001
MM202 21 106 466 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=12219  $PIN_XY=13134,12222,13104,12219,13074,12222 $DEVICE_ID=1001
MM203 GND! 412 231 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=11844  $PIN_XY=13134,11928,13104,11844,13074,11928 $DEVICE_ID=1001
MM204 21 105 412 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=11295  $PIN_XY=13134,11298,13104,11295,13074,11298 $DEVICE_ID=1001
MM205 GND! 417 236 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=10920  $PIN_XY=13134,11004,13104,10920,13074,11004 $DEVICE_ID=1001
MM206 21 104 417 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=10371  $PIN_XY=13134,10374,13104,10371,13074,10374 $DEVICE_ID=1001
MM207 GND! 420 160 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=9996  $PIN_XY=13134,10080,13104,9996,13074,10080 $DEVICE_ID=1001
MM208 21 103 420 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=9447  $PIN_XY=13134,9450,13104,9447,13074,9450 $DEVICE_ID=1001
MM209 GND! 366 159 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=9072  $PIN_XY=13134,9156,13104,9072,13074,9156 $DEVICE_ID=1001
MM210 21 99 366 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=8523  $PIN_XY=13134,8526,13104,8523,13074,8526 $DEVICE_ID=1001
MM211 224 108 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=14703  $PIN_XY=12966,14700,12936,14703,12906,14700 $DEVICE_ID=1001
MM212 462 224 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=14154  $PIN_XY=12966,14070,12936,14154,12906,14070 $DEVICE_ID=1001
MM213 227 107 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=13779  $PIN_XY=12966,13776,12936,13779,12906,13776 $DEVICE_ID=1001
MM214 465 227 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=13230  $PIN_XY=12966,13146,12936,13230,12906,13146 $DEVICE_ID=1001
MM215 228 106 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=12855  $PIN_XY=12966,12852,12936,12855,12906,12852 $DEVICE_ID=1001
MM216 466 228 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=12306  $PIN_XY=12966,12222,12936,12306,12906,12222 $DEVICE_ID=1001
MM217 231 105 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=11931  $PIN_XY=12966,11928,12936,11931,12906,11928 $DEVICE_ID=1001
MM218 412 231 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=11382  $PIN_XY=12966,11298,12936,11382,12906,11298 $DEVICE_ID=1001
MM219 236 104 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=11007  $PIN_XY=12966,11004,12936,11007,12906,11004 $DEVICE_ID=1001
MM220 417 236 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=10458  $PIN_XY=12966,10374,12936,10458,12906,10374 $DEVICE_ID=1001
MM221 160 103 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=10083  $PIN_XY=12966,10080,12936,10083,12906,10080 $DEVICE_ID=1001
MM222 420 160 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=9534  $PIN_XY=12966,9450,12936,9534,12906,9450 $DEVICE_ID=1001
MM223 159 99 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=9159  $PIN_XY=12966,9156,12936,9159,12906,9156 $DEVICE_ID=1001
MM224 366 159 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=8610  $PIN_XY=12966,8526,12936,8610,12906,8526 $DEVICE_ID=1001
MM225 GND! 435 199 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=14616  $PIN_XY=12126,14700,12096,14616,12066,14700 $DEVICE_ID=1001
MM226 17 108 435 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=14067  $PIN_XY=12126,14070,12096,14067,12066,14070 $DEVICE_ID=1001
MM227 GND! 437 201 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=13692  $PIN_XY=12126,13776,12096,13692,12066,13776 $DEVICE_ID=1001
MM228 17 107 437 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=13143  $PIN_XY=12126,13146,12096,13143,12066,13146 $DEVICE_ID=1001
MM229 GND! 442 206 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=12768  $PIN_XY=12126,12852,12096,12768,12066,12852 $DEVICE_ID=1001
MM230 17 106 442 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=12219  $PIN_XY=12126,12222,12096,12219,12066,12222 $DEVICE_ID=1001
MM231 GND! 388 212 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=11844  $PIN_XY=12126,11928,12096,11844,12066,11928 $DEVICE_ID=1001
MM232 199 108 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=14703  $PIN_XY=11958,14700,11928,14703,11898,14700 $DEVICE_ID=1001
MM233 435 199 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=14154  $PIN_XY=11958,14070,11928,14154,11898,14070 $DEVICE_ID=1001
MM234 201 107 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=13779  $PIN_XY=11958,13776,11928,13779,11898,13776 $DEVICE_ID=1001
MM235 437 201 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=13230  $PIN_XY=11958,13146,11928,13230,11898,13146 $DEVICE_ID=1001
MM236 206 106 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=12855  $PIN_XY=11958,12852,11928,12855,11898,12852 $DEVICE_ID=1001
MM237 442 206 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=12306  $PIN_XY=11958,12222,11928,12306,11898,12222 $DEVICE_ID=1001
MM238 212 105 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=11931  $PIN_XY=11958,11928,11928,11931,11898,11928 $DEVICE_ID=1001
MM239 GND! 434 198 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=14616  $PIN_XY=11454,14700,11424,14616,11394,14700 $DEVICE_ID=1001
MM240 16 108 434 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=14067  $PIN_XY=11454,14070,11424,14067,11394,14070 $DEVICE_ID=1001
MM241 GND! 438 202 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=13692  $PIN_XY=11454,13776,11424,13692,11394,13776 $DEVICE_ID=1001
MM242 16 107 438 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=13143  $PIN_XY=11454,13146,11424,13143,11394,13146 $DEVICE_ID=1001
MM243 GND! 443 207 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=12768  $PIN_XY=11454,12852,11424,12768,11394,12852 $DEVICE_ID=1001
MM244 16 106 443 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=12219  $PIN_XY=11454,12222,11424,12219,11394,12222 $DEVICE_ID=1001
MM245 GND! 387 211 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=11844  $PIN_XY=11454,11928,11424,11844,11394,11928 $DEVICE_ID=1001
MM246 198 108 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=14703  $PIN_XY=11286,14700,11256,14703,11226,14700 $DEVICE_ID=1001
MM247 434 198 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=14154  $PIN_XY=11286,14070,11256,14154,11226,14070 $DEVICE_ID=1001
MM248 202 107 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=13779  $PIN_XY=11286,13776,11256,13779,11226,13776 $DEVICE_ID=1001
MM249 438 202 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=13230  $PIN_XY=11286,13146,11256,13230,11226,13146 $DEVICE_ID=1001
MM250 207 106 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=12855  $PIN_XY=11286,12852,11256,12855,11226,12852 $DEVICE_ID=1001
MM251 443 207 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=12306  $PIN_XY=11286,12222,11256,12306,11226,12222 $DEVICE_ID=1001
MM252 211 105 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=11931  $PIN_XY=11286,11928,11256,11931,11226,11928 $DEVICE_ID=1001
MM253 GND! 433 197 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=14616  $PIN_XY=10782,14700,10752,14616,10722,14700 $DEVICE_ID=1001
MM254 15 108 433 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=14067  $PIN_XY=10782,14070,10752,14067,10722,14070 $DEVICE_ID=1001
MM255 GND! 439 203 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=13692  $PIN_XY=10782,13776,10752,13692,10722,13776 $DEVICE_ID=1001
MM256 15 107 439 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=13143  $PIN_XY=10782,13146,10752,13143,10722,13146 $DEVICE_ID=1001
MM257 GND! 444 208 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=12768  $PIN_XY=10782,12852,10752,12768,10722,12852 $DEVICE_ID=1001
MM258 15 106 444 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=12219  $PIN_XY=10782,12222,10752,12219,10722,12222 $DEVICE_ID=1001
MM259 GND! 386 210 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=11844  $PIN_XY=10782,11928,10752,11844,10722,11928 $DEVICE_ID=1001
MM260 197 108 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=14703  $PIN_XY=10614,14700,10584,14703,10554,14700 $DEVICE_ID=1001
MM261 433 197 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=14154  $PIN_XY=10614,14070,10584,14154,10554,14070 $DEVICE_ID=1001
MM262 203 107 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=13779  $PIN_XY=10614,13776,10584,13779,10554,13776 $DEVICE_ID=1001
MM263 439 203 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=13230  $PIN_XY=10614,13146,10584,13230,10554,13146 $DEVICE_ID=1001
MM264 208 106 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=12855  $PIN_XY=10614,12852,10584,12855,10554,12852 $DEVICE_ID=1001
MM265 444 208 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=12306  $PIN_XY=10614,12222,10584,12306,10554,12222 $DEVICE_ID=1001
MM266 210 105 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=11931  $PIN_XY=10614,11928,10584,11931,10554,11928 $DEVICE_ID=1001
MM267 17 105 388 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=11295  $PIN_XY=12126,11298,12096,11295,12066,11298 $DEVICE_ID=1001
MM268 GND! 391 215 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=10920  $PIN_XY=12126,11004,12096,10920,12066,11004 $DEVICE_ID=1001
MM269 17 104 391 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=10371  $PIN_XY=12126,10374,12096,10371,12066,10374 $DEVICE_ID=1001
MM270 GND! 393 152 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=9996  $PIN_XY=12126,10080,12096,9996,12066,10080 $DEVICE_ID=1001
MM271 17 103 393 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=9447  $PIN_XY=12126,9450,12096,9447,12066,9450 $DEVICE_ID=1001
MM272 GND! 352 151 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=9072  $PIN_XY=12126,9156,12096,9072,12066,9156 $DEVICE_ID=1001
MM273 17 99 352 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=8523  $PIN_XY=12126,8526,12096,8523,12066,8526 $DEVICE_ID=1001
MM274 388 212 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=11382  $PIN_XY=11958,11298,11928,11382,11898,11298 $DEVICE_ID=1001
MM275 215 104 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=11007  $PIN_XY=11958,11004,11928,11007,11898,11004 $DEVICE_ID=1001
MM276 391 215 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=10458  $PIN_XY=11958,10374,11928,10458,11898,10374 $DEVICE_ID=1001
MM277 152 103 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=10083  $PIN_XY=11958,10080,11928,10083,11898,10080 $DEVICE_ID=1001
MM278 393 152 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=9534  $PIN_XY=11958,9450,11928,9534,11898,9450 $DEVICE_ID=1001
MM279 151 99 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=9159  $PIN_XY=11958,9156,11928,9159,11898,9156 $DEVICE_ID=1001
MM280 352 151 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=8610  $PIN_XY=11958,8526,11928,8610,11898,8526 $DEVICE_ID=1001
MM281 16 105 387 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=11295  $PIN_XY=11454,11298,11424,11295,11394,11298 $DEVICE_ID=1001
MM282 GND! 390 214 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=10920  $PIN_XY=11454,11004,11424,10920,11394,11004 $DEVICE_ID=1001
MM283 16 104 390 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=10371  $PIN_XY=11454,10374,11424,10371,11394,10374 $DEVICE_ID=1001
MM284 GND! 394 150 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=9996  $PIN_XY=11454,10080,11424,9996,11394,10080 $DEVICE_ID=1001
MM285 16 103 394 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=9447  $PIN_XY=11454,9450,11424,9447,11394,9450 $DEVICE_ID=1001
MM286 GND! 351 149 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=9072  $PIN_XY=11454,9156,11424,9072,11394,9156 $DEVICE_ID=1001
MM287 16 99 351 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=8523  $PIN_XY=11454,8526,11424,8523,11394,8526 $DEVICE_ID=1001
MM288 387 211 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=11382  $PIN_XY=11286,11298,11256,11382,11226,11298 $DEVICE_ID=1001
MM289 214 104 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=11007  $PIN_XY=11286,11004,11256,11007,11226,11004 $DEVICE_ID=1001
MM290 390 214 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=10458  $PIN_XY=11286,10374,11256,10458,11226,10374 $DEVICE_ID=1001
MM291 150 103 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=10083  $PIN_XY=11286,10080,11256,10083,11226,10080 $DEVICE_ID=1001
MM292 394 150 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=9534  $PIN_XY=11286,9450,11256,9534,11226,9450 $DEVICE_ID=1001
MM293 149 99 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=9159  $PIN_XY=11286,9156,11256,9159,11226,9156 $DEVICE_ID=1001
MM294 351 149 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=8610  $PIN_XY=11286,8526,11256,8610,11226,8526 $DEVICE_ID=1001
MM295 15 105 386 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=11295  $PIN_XY=10782,11298,10752,11295,10722,11298 $DEVICE_ID=1001
MM296 GND! 389 213 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=10920  $PIN_XY=10782,11004,10752,10920,10722,11004 $DEVICE_ID=1001
MM297 15 104 389 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=10371  $PIN_XY=10782,10374,10752,10371,10722,10374 $DEVICE_ID=1001
MM298 GND! 395 148 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=9996  $PIN_XY=10782,10080,10752,9996,10722,10080 $DEVICE_ID=1001
MM299 15 103 395 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=9447  $PIN_XY=10782,9450,10752,9447,10722,9450 $DEVICE_ID=1001
MM300 GND! 350 147 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=9072  $PIN_XY=10782,9156,10752,9072,10722,9156 $DEVICE_ID=1001
MM301 15 99 350 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=8523  $PIN_XY=10782,8526,10752,8523,10722,8526 $DEVICE_ID=1001
MM302 386 210 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=11382  $PIN_XY=10614,11298,10584,11382,10554,11298 $DEVICE_ID=1001
MM303 213 104 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=11007  $PIN_XY=10614,11004,10584,11007,10554,11004 $DEVICE_ID=1001
MM304 389 213 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=10458  $PIN_XY=10614,10374,10584,10458,10554,10374 $DEVICE_ID=1001
MM305 148 103 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=10083  $PIN_XY=10614,10080,10584,10083,10554,10080 $DEVICE_ID=1001
MM306 395 148 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=9534  $PIN_XY=10614,9450,10584,9534,10554,9450 $DEVICE_ID=1001
MM307 147 99 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=9159  $PIN_XY=10614,9156,10584,9159,10554,9156 $DEVICE_ID=1001
MM308 350 147 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=8610  $PIN_XY=10614,8526,10584,8610,10554,8526 $DEVICE_ID=1001
MM309 GND! 436 200 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=14616  $PIN_XY=10110,14700,10080,14616,10050,14700 $DEVICE_ID=1001
MM310 13 108 436 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=14067  $PIN_XY=10110,14070,10080,14067,10050,14070 $DEVICE_ID=1001
MM311 GND! 440 204 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=13692  $PIN_XY=10110,13776,10080,13692,10050,13776 $DEVICE_ID=1001
MM312 13 107 440 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=13143  $PIN_XY=10110,13146,10080,13143,10050,13146 $DEVICE_ID=1001
MM313 GND! 441 205 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=12768  $PIN_XY=10110,12852,10080,12768,10050,12852 $DEVICE_ID=1001
MM314 13 106 441 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=12219  $PIN_XY=10110,12222,10080,12219,10050,12222 $DEVICE_ID=1001
MM315 GND! 385 209 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=11844  $PIN_XY=10110,11928,10080,11844,10050,11928 $DEVICE_ID=1001
MM316 200 108 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=14703  $PIN_XY=9942,14700,9912,14703,9882,14700 $DEVICE_ID=1001
MM317 436 200 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=14154  $PIN_XY=9942,14070,9912,14154,9882,14070 $DEVICE_ID=1001
MM318 204 107 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=13779  $PIN_XY=9942,13776,9912,13779,9882,13776 $DEVICE_ID=1001
MM319 440 204 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=13230  $PIN_XY=9942,13146,9912,13230,9882,13146 $DEVICE_ID=1001
MM320 205 106 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=12855  $PIN_XY=9942,12852,9912,12855,9882,12852 $DEVICE_ID=1001
MM321 441 205 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=12306  $PIN_XY=9942,12222,9912,12306,9882,12222 $DEVICE_ID=1001
MM322 209 105 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=11931  $PIN_XY=9942,11928,9912,11931,9882,11928 $DEVICE_ID=1001
MM323 GND! 430 196 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=14616  $PIN_XY=9102,14700,9072,14616,9042,14700 $DEVICE_ID=1001
MM324 8 108 430 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=14067  $PIN_XY=9102,14070,9072,14067,9042,14070 $DEVICE_ID=1001
MM325 GND! 428 191 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=13692  $PIN_XY=9102,13776,9072,13692,9042,13776 $DEVICE_ID=1001
MM326 8 107 428 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=13143  $PIN_XY=9102,13146,9072,13143,9042,13146 $DEVICE_ID=1001
MM327 GND! 423 185 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=12768  $PIN_XY=9102,12852,9072,12768,9042,12852 $DEVICE_ID=1001
MM328 8 106 423 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=12219  $PIN_XY=9102,12222,9072,12219,9042,12222 $DEVICE_ID=1001
MM329 GND! 381 182 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=11844  $PIN_XY=9102,11928,9072,11844,9042,11928 $DEVICE_ID=1001
MM330 196 108 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=14703  $PIN_XY=8934,14700,8904,14703,8874,14700 $DEVICE_ID=1001
MM331 430 196 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=14154  $PIN_XY=8934,14070,8904,14154,8874,14070 $DEVICE_ID=1001
MM332 191 107 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=13779  $PIN_XY=8934,13776,8904,13779,8874,13776 $DEVICE_ID=1001
MM333 428 191 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=13230  $PIN_XY=8934,13146,8904,13230,8874,13146 $DEVICE_ID=1001
MM334 185 106 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=12855  $PIN_XY=8934,12852,8904,12855,8874,12852 $DEVICE_ID=1001
MM335 423 185 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=12306  $PIN_XY=8934,12222,8904,12306,8874,12222 $DEVICE_ID=1001
MM336 182 105 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=11931  $PIN_XY=8934,11928,8904,11931,8874,11928 $DEVICE_ID=1001
MM337 GND! 431 195 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=14616  $PIN_XY=8430,14700,8400,14616,8370,14700 $DEVICE_ID=1001
MM338 10 108 431 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=14067  $PIN_XY=8430,14070,8400,14067,8370,14070 $DEVICE_ID=1001
MM339 GND! 427 190 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=13692  $PIN_XY=8430,13776,8400,13692,8370,13776 $DEVICE_ID=1001
MM340 10 107 427 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=13143  $PIN_XY=8430,13146,8400,13143,8370,13146 $DEVICE_ID=1001
MM341 GND! 422 186 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=12768  $PIN_XY=8430,12852,8400,12768,8370,12852 $DEVICE_ID=1001
MM342 10 106 422 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=12219  $PIN_XY=8430,12222,8400,12219,8370,12222 $DEVICE_ID=1001
MM343 GND! 382 183 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=11844  $PIN_XY=8430,11928,8400,11844,8370,11928 $DEVICE_ID=1001
MM344 13 105 385 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=11295  $PIN_XY=10110,11298,10080,11295,10050,11298 $DEVICE_ID=1001
MM345 GND! 392 216 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=10920  $PIN_XY=10110,11004,10080,10920,10050,11004 $DEVICE_ID=1001
MM346 13 104 392 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=10371  $PIN_XY=10110,10374,10080,10371,10050,10374 $DEVICE_ID=1001
MM347 GND! 396 146 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=9996  $PIN_XY=10110,10080,10080,9996,10050,10080 $DEVICE_ID=1001
MM348 13 103 396 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=9447  $PIN_XY=10110,9450,10080,9447,10050,9450 $DEVICE_ID=1001
MM349 GND! 349 145 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=9072  $PIN_XY=10110,9156,10080,9072,10050,9156 $DEVICE_ID=1001
MM350 13 99 349 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=8523  $PIN_XY=10110,8526,10080,8523,10050,8526 $DEVICE_ID=1001
MM351 385 209 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=11382  $PIN_XY=9942,11298,9912,11382,9882,11298 $DEVICE_ID=1001
MM352 216 104 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=11007  $PIN_XY=9942,11004,9912,11007,9882,11004 $DEVICE_ID=1001
MM353 392 216 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=10458  $PIN_XY=9942,10374,9912,10458,9882,10374 $DEVICE_ID=1001
MM354 146 103 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=10083  $PIN_XY=9942,10080,9912,10083,9882,10080 $DEVICE_ID=1001
MM355 396 146 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=9534  $PIN_XY=9942,9450,9912,9534,9882,9450 $DEVICE_ID=1001
MM356 145 99 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=9159  $PIN_XY=9942,9156,9912,9159,9882,9156 $DEVICE_ID=1001
MM357 349 145 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=8610  $PIN_XY=9942,8526,9912,8610,9882,8526 $DEVICE_ID=1001
MM358 8 105 381 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=11295  $PIN_XY=9102,11298,9072,11295,9042,11298 $DEVICE_ID=1001
MM359 GND! 378 180 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=10920  $PIN_XY=9102,11004,9072,10920,9042,11004 $DEVICE_ID=1001
MM360 8 104 378 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=10371  $PIN_XY=9102,10374,9072,10371,9042,10374 $DEVICE_ID=1001
MM361 GND! 376 138 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=9996  $PIN_XY=9102,10080,9072,9996,9042,10080 $DEVICE_ID=1001
MM362 8 103 376 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=9447  $PIN_XY=9102,9450,9072,9447,9042,9450 $DEVICE_ID=1001
MM363 GND! 346 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=9072  $PIN_XY=9102,9156,9072,9072,9042,9156 $DEVICE_ID=1001
MM364 8 99 346 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=8523  $PIN_XY=9102,8526,9072,8523,9042,8526 $DEVICE_ID=1001
MM365 381 182 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=11382  $PIN_XY=8934,11298,8904,11382,8874,11298 $DEVICE_ID=1001
MM366 180 104 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=11007  $PIN_XY=8934,11004,8904,11007,8874,11004 $DEVICE_ID=1001
MM367 378 180 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=10458  $PIN_XY=8934,10374,8904,10458,8874,10374 $DEVICE_ID=1001
MM368 138 103 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=10083  $PIN_XY=8934,10080,8904,10083,8874,10080 $DEVICE_ID=1001
MM369 376 138 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=9534  $PIN_XY=8934,9450,8904,9534,8874,9450 $DEVICE_ID=1001
MM370 133 99 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=9159  $PIN_XY=8934,9156,8904,9159,8874,9156 $DEVICE_ID=1001
MM371 346 133 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=8610  $PIN_XY=8934,8526,8904,8610,8874,8526 $DEVICE_ID=1001
MM372 10 105 382 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=11295  $PIN_XY=8430,11298,8400,11295,8370,11298 $DEVICE_ID=1001
MM373 GND! 379 179 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=10920  $PIN_XY=8430,11004,8400,10920,8370,11004 $DEVICE_ID=1001
MM374 10 104 379 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=10371  $PIN_XY=8430,10374,8400,10371,8370,10374 $DEVICE_ID=1001
MM375 GND! 375 137 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=9996  $PIN_XY=8430,10080,8400,9996,8370,10080 $DEVICE_ID=1001
MM376 10 103 375 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=9447  $PIN_XY=8430,9450,8400,9447,8370,9450 $DEVICE_ID=1001
MM377 GND! 345 134 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=9072  $PIN_XY=8430,9156,8400,9072,8370,9156 $DEVICE_ID=1001
MM378 10 99 345 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=8523  $PIN_XY=8430,8526,8400,8523,8370,8526 $DEVICE_ID=1001
MM379 195 108 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=14703  $PIN_XY=8262,14700,8232,14703,8202,14700 $DEVICE_ID=1001
MM380 431 195 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=14154  $PIN_XY=8262,14070,8232,14154,8202,14070 $DEVICE_ID=1001
MM381 190 107 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=13779  $PIN_XY=8262,13776,8232,13779,8202,13776 $DEVICE_ID=1001
MM382 427 190 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=13230  $PIN_XY=8262,13146,8232,13230,8202,13146 $DEVICE_ID=1001
MM383 186 106 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=12855  $PIN_XY=8262,12852,8232,12855,8202,12852 $DEVICE_ID=1001
MM384 422 186 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=12306  $PIN_XY=8262,12222,8232,12306,8202,12222 $DEVICE_ID=1001
MM385 183 105 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=11931  $PIN_XY=8262,11928,8232,11931,8202,11928 $DEVICE_ID=1001
MM386 GND! 432 194 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=14616  $PIN_XY=7758,14700,7728,14616,7698,14700 $DEVICE_ID=1001
MM387 11 108 432 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=14067  $PIN_XY=7758,14070,7728,14067,7698,14070 $DEVICE_ID=1001
MM388 GND! 426 189 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=13692  $PIN_XY=7758,13776,7728,13692,7698,13776 $DEVICE_ID=1001
MM389 11 107 426 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=13143  $PIN_XY=7758,13146,7728,13143,7698,13146 $DEVICE_ID=1001
MM390 GND! 421 187 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=12768  $PIN_XY=7758,12852,7728,12768,7698,12852 $DEVICE_ID=1001
MM391 11 106 421 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=12219  $PIN_XY=7758,12222,7728,12219,7698,12222 $DEVICE_ID=1001
MM392 GND! 383 184 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=11844  $PIN_XY=7758,11928,7728,11844,7698,11928 $DEVICE_ID=1001
MM393 194 108 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=14703  $PIN_XY=7590,14700,7560,14703,7530,14700 $DEVICE_ID=1001
MM394 432 194 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=14154  $PIN_XY=7590,14070,7560,14154,7530,14070 $DEVICE_ID=1001
MM395 189 107 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=13779  $PIN_XY=7590,13776,7560,13779,7530,13776 $DEVICE_ID=1001
MM396 426 189 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=13230  $PIN_XY=7590,13146,7560,13230,7530,13146 $DEVICE_ID=1001
MM397 187 106 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=12855  $PIN_XY=7590,12852,7560,12855,7530,12852 $DEVICE_ID=1001
MM398 421 187 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=12306  $PIN_XY=7590,12222,7560,12306,7530,12222 $DEVICE_ID=1001
MM399 184 105 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=11931  $PIN_XY=7590,11928,7560,11931,7530,11928 $DEVICE_ID=1001
MM400 GND! 429 193 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=14616  $PIN_XY=7086,14700,7056,14616,7026,14700 $DEVICE_ID=1001
MM401 12 108 429 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=14067  $PIN_XY=7086,14070,7056,14067,7026,14070 $DEVICE_ID=1001
MM402 GND! 425 192 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=13692  $PIN_XY=7086,13776,7056,13692,7026,13776 $DEVICE_ID=1001
MM403 12 107 425 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=13143  $PIN_XY=7086,13146,7056,13143,7026,13146 $DEVICE_ID=1001
MM404 GND! 424 188 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=12768  $PIN_XY=7086,12852,7056,12768,7026,12852 $DEVICE_ID=1001
MM405 12 106 424 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=12219  $PIN_XY=7086,12222,7056,12219,7026,12222 $DEVICE_ID=1001
MM406 GND! 384 181 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=11844  $PIN_XY=7086,11928,7056,11844,7026,11928 $DEVICE_ID=1001
MM407 193 108 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=14703  $PIN_XY=6918,14700,6888,14703,6858,14700 $DEVICE_ID=1001
MM408 429 193 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=14154  $PIN_XY=6918,14070,6888,14154,6858,14070 $DEVICE_ID=1001
MM409 192 107 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=13779  $PIN_XY=6918,13776,6888,13779,6858,13776 $DEVICE_ID=1001
MM410 425 192 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=13230  $PIN_XY=6918,13146,6888,13230,6858,13146 $DEVICE_ID=1001
MM411 188 106 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=12855  $PIN_XY=6918,12852,6888,12855,6858,12852 $DEVICE_ID=1001
MM412 424 188 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=12306  $PIN_XY=6918,12222,6888,12306,6858,12222 $DEVICE_ID=1001
MM413 181 105 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=11931  $PIN_XY=6918,11928,6888,11931,6858,11928 $DEVICE_ID=1001
MM414 382 183 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=11382  $PIN_XY=8262,11298,8232,11382,8202,11298 $DEVICE_ID=1001
MM415 179 104 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=11007  $PIN_XY=8262,11004,8232,11007,8202,11004 $DEVICE_ID=1001
MM416 379 179 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=10458  $PIN_XY=8262,10374,8232,10458,8202,10374 $DEVICE_ID=1001
MM417 137 103 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=10083  $PIN_XY=8262,10080,8232,10083,8202,10080 $DEVICE_ID=1001
MM418 375 137 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=9534  $PIN_XY=8262,9450,8232,9534,8202,9450 $DEVICE_ID=1001
MM419 134 99 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=9159  $PIN_XY=8262,9156,8232,9159,8202,9156 $DEVICE_ID=1001
MM420 345 134 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=8610  $PIN_XY=8262,8526,8232,8610,8202,8526 $DEVICE_ID=1001
MM421 11 105 383 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=11295  $PIN_XY=7758,11298,7728,11295,7698,11298 $DEVICE_ID=1001
MM422 GND! 380 178 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=10920  $PIN_XY=7758,11004,7728,10920,7698,11004 $DEVICE_ID=1001
MM423 11 104 380 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=10371  $PIN_XY=7758,10374,7728,10371,7698,10374 $DEVICE_ID=1001
MM424 GND! 374 136 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=9996  $PIN_XY=7758,10080,7728,9996,7698,10080 $DEVICE_ID=1001
MM425 11 103 374 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=9447  $PIN_XY=7758,9450,7728,9447,7698,9450 $DEVICE_ID=1001
MM426 GND! 344 135 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=9072  $PIN_XY=7758,9156,7728,9072,7698,9156 $DEVICE_ID=1001
MM427 11 99 344 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=8523  $PIN_XY=7758,8526,7728,8523,7698,8526 $DEVICE_ID=1001
MM428 383 184 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=11382  $PIN_XY=7590,11298,7560,11382,7530,11298 $DEVICE_ID=1001
MM429 178 104 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=11007  $PIN_XY=7590,11004,7560,11007,7530,11004 $DEVICE_ID=1001
MM430 380 178 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=10458  $PIN_XY=7590,10374,7560,10458,7530,10374 $DEVICE_ID=1001
MM431 136 103 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=10083  $PIN_XY=7590,10080,7560,10083,7530,10080 $DEVICE_ID=1001
MM432 374 136 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=9534  $PIN_XY=7590,9450,7560,9534,7530,9450 $DEVICE_ID=1001
MM433 135 99 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=9159  $PIN_XY=7590,9156,7560,9159,7530,9156 $DEVICE_ID=1001
MM434 344 135 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=8610  $PIN_XY=7590,8526,7560,8610,7530,8526 $DEVICE_ID=1001
MM435 12 105 384 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=11295  $PIN_XY=7086,11298,7056,11295,7026,11298 $DEVICE_ID=1001
MM436 GND! 377 177 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=10920  $PIN_XY=7086,11004,7056,10920,7026,11004 $DEVICE_ID=1001
MM437 12 104 377 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=10371  $PIN_XY=7086,10374,7056,10371,7026,10374 $DEVICE_ID=1001
MM438 GND! 373 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=9996  $PIN_XY=7086,10080,7056,9996,7026,10080 $DEVICE_ID=1001
MM439 12 103 373 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=9447  $PIN_XY=7086,9450,7056,9447,7026,9450 $DEVICE_ID=1001
MM440 GND! 348 139 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=9072  $PIN_XY=7086,9156,7056,9072,7026,9156 $DEVICE_ID=1001
MM441 12 99 348 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=8523  $PIN_XY=7086,8526,7056,8523,7026,8526 $DEVICE_ID=1001
MM442 384 181 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=11382  $PIN_XY=6918,11298,6888,11382,6858,11298 $DEVICE_ID=1001
MM443 177 104 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=11007  $PIN_XY=6918,11004,6888,11007,6858,11004 $DEVICE_ID=1001
MM444 377 177 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=10458  $PIN_XY=6918,10374,6888,10458,6858,10374 $DEVICE_ID=1001
MM445 140 103 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=10083  $PIN_XY=6918,10080,6888,10083,6858,10080 $DEVICE_ID=1001
MM446 373 140 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=9534  $PIN_XY=6918,9450,6888,9534,6858,9450 $DEVICE_ID=1001
MM447 139 99 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=9159  $PIN_XY=6918,9156,6888,9159,6858,9156 $DEVICE_ID=1001
MM448 348 139 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=8610  $PIN_XY=6918,8526,6888,8610,6858,8526 $DEVICE_ID=1001
MM449 GND! 365 500 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=8148  $PIN_XY=18174,8232,18144,8148,18114,8232 $DEVICE_ID=1001
MM450 27 98 365 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=7620  $PIN_XY=18174,7602,18144,7620,18114,7602 $DEVICE_ID=1001
MM451 500 98 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=8235  $PIN_XY=18006,8232,17976,8235,17946,8232 $DEVICE_ID=1001
MM452 365 500 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=7707  $PIN_XY=18006,7602,17976,7707,17946,7602 $DEVICE_ID=1001
MM453 GND! 364 499 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=8148  $PIN_XY=17502,8232,17472,8148,17442,8232 $DEVICE_ID=1001
MM454 26 98 364 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=7620  $PIN_XY=17502,7602,17472,7620,17442,7602 $DEVICE_ID=1001
MM455 499 98 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=8235  $PIN_XY=17334,8232,17304,8235,17274,8232 $DEVICE_ID=1001
MM456 364 499 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=7707  $PIN_XY=17334,7602,17304,7707,17274,7602 $DEVICE_ID=1001
MM457 GND! 363 498 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=8148  $PIN_XY=16830,8232,16800,8148,16770,8232 $DEVICE_ID=1001
MM458 25 98 363 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=7620  $PIN_XY=16830,7602,16800,7620,16770,7602 $DEVICE_ID=1001
MM459 498 98 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=8235  $PIN_XY=16662,8232,16632,8235,16602,8232 $DEVICE_ID=1001
MM460 363 498 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=7707  $PIN_XY=16662,7602,16632,7707,16602,7602 $DEVICE_ID=1001
MM461 GND! 362 497 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=8148  $PIN_XY=16158,8232,16128,8148,16098,8232 $DEVICE_ID=1001
MM462 23 98 362 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=7620  $PIN_XY=16158,7602,16128,7620,16098,7602 $DEVICE_ID=1001
MM463 497 98 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=8235  $PIN_XY=15990,8232,15960,8235,15930,8232 $DEVICE_ID=1001
MM464 362 497 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=7707  $PIN_XY=15990,7602,15960,7707,15930,7602 $DEVICE_ID=1001
MM465 GND! 369 501 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=8148  $PIN_XY=15150,8232,15120,8148,15090,8232 $DEVICE_ID=1001
MM466 22 98 369 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=7620  $PIN_XY=15150,7602,15120,7620,15090,7602 $DEVICE_ID=1001
MM467 501 98 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=8235  $PIN_XY=14982,8232,14952,8235,14922,8232 $DEVICE_ID=1001
MM468 369 501 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=7707  $PIN_XY=14982,7602,14952,7707,14922,7602 $DEVICE_ID=1001
MM469 GND! 370 502 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=8148  $PIN_XY=14478,8232,14448,8148,14418,8232 $DEVICE_ID=1001
MM470 18 98 370 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=7620  $PIN_XY=14478,7602,14448,7620,14418,7602 $DEVICE_ID=1001
MM471 502 98 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=8235  $PIN_XY=14310,8232,14280,8235,14250,8232 $DEVICE_ID=1001
MM472 370 502 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=7707  $PIN_XY=14310,7602,14280,7707,14250,7602 $DEVICE_ID=1001
MM473 GND! 371 495 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=8148  $PIN_XY=13806,8232,13776,8148,13746,8232 $DEVICE_ID=1001
MM474 20 98 371 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=7620  $PIN_XY=13806,7602,13776,7620,13746,7602 $DEVICE_ID=1001
MM475 495 98 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=8235  $PIN_XY=13638,8232,13608,8235,13578,8232 $DEVICE_ID=1001
MM476 371 495 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=7707  $PIN_XY=13638,7602,13608,7707,13578,7602 $DEVICE_ID=1001
MM477 GND! 372 496 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=8148  $PIN_XY=13134,8232,13104,8148,13074,8232 $DEVICE_ID=1001
MM478 21 98 372 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=7620  $PIN_XY=13134,7602,13104,7620,13074,7602 $DEVICE_ID=1001
MM479 496 98 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=8235  $PIN_XY=12966,8232,12936,8235,12906,8232 $DEVICE_ID=1001
MM480 372 496 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=7707  $PIN_XY=12966,7602,12936,7707,12906,7602 $DEVICE_ID=1001
MM481 GND! 353 491 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=8148  $PIN_XY=12126,8232,12096,8148,12066,8232 $DEVICE_ID=1001
MM482 17 98 353 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=7620  $PIN_XY=12126,7602,12096,7620,12066,7602 $DEVICE_ID=1001
MM483 491 98 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=8235  $PIN_XY=11958,8232,11928,8235,11898,8232 $DEVICE_ID=1001
MM484 353 491 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=7707  $PIN_XY=11958,7602,11928,7707,11898,7602 $DEVICE_ID=1001
MM485 GND! 354 492 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=8148  $PIN_XY=11454,8232,11424,8148,11394,8232 $DEVICE_ID=1001
MM486 16 98 354 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=7620  $PIN_XY=11454,7602,11424,7620,11394,7602 $DEVICE_ID=1001
MM487 492 98 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=8235  $PIN_XY=11286,8232,11256,8235,11226,8232 $DEVICE_ID=1001
MM488 354 492 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=7707  $PIN_XY=11286,7602,11256,7707,11226,7602 $DEVICE_ID=1001
MM489 GND! 355 493 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=8148  $PIN_XY=10782,8232,10752,8148,10722,8232 $DEVICE_ID=1001
MM490 15 98 355 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=7620  $PIN_XY=10782,7602,10752,7620,10722,7602 $DEVICE_ID=1001
MM491 493 98 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=8235  $PIN_XY=10614,8232,10584,8235,10554,8232 $DEVICE_ID=1001
MM492 355 493 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=7707  $PIN_XY=10614,7602,10584,7707,10554,7602 $DEVICE_ID=1001
MM493 GND! 356 494 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=8148  $PIN_XY=10110,8232,10080,8148,10050,8232 $DEVICE_ID=1001
MM494 13 98 356 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=7620  $PIN_XY=10110,7602,10080,7620,10050,7602 $DEVICE_ID=1001
MM495 494 98 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=8235  $PIN_XY=9942,8232,9912,8235,9882,8232 $DEVICE_ID=1001
MM496 356 494 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=7707  $PIN_XY=9942,7602,9912,7707,9882,7602 $DEVICE_ID=1001
MM497 GND! 341 487 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=8148  $PIN_XY=9102,8232,9072,8148,9042,8232 $DEVICE_ID=1001
MM498 8 98 341 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=7620  $PIN_XY=9102,7602,9072,7620,9042,7602 $DEVICE_ID=1001
MM499 487 98 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=8235  $PIN_XY=8934,8232,8904,8235,8874,8232 $DEVICE_ID=1001
MM500 341 487 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=7707  $PIN_XY=8934,7602,8904,7707,8874,7602 $DEVICE_ID=1001
MM501 GND! 342 488 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=8148  $PIN_XY=8430,8232,8400,8148,8370,8232 $DEVICE_ID=1001
MM502 10 98 342 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=7620  $PIN_XY=8430,7602,8400,7620,8370,7602 $DEVICE_ID=1001
MM503 488 98 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=8235  $PIN_XY=8262,8232,8232,8235,8202,8232 $DEVICE_ID=1001
MM504 342 488 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=7707  $PIN_XY=8262,7602,8232,7707,8202,7602 $DEVICE_ID=1001
MM505 GND! 343 489 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=8148  $PIN_XY=7758,8232,7728,8148,7698,8232 $DEVICE_ID=1001
MM506 11 98 343 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=7620  $PIN_XY=7758,7602,7728,7620,7698,7602 $DEVICE_ID=1001
MM507 489 98 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=8235  $PIN_XY=7590,8232,7560,8235,7530,8232 $DEVICE_ID=1001
MM508 343 489 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=7707  $PIN_XY=7590,7602,7560,7707,7530,7602 $DEVICE_ID=1001
MM509 GND! 347 490 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=8148  $PIN_XY=7086,8232,7056,8148,7026,8232 $DEVICE_ID=1001
MM510 12 98 347 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=7620  $PIN_XY=7086,7602,7056,7620,7026,7602 $DEVICE_ID=1001
MM511 490 98 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=8235  $PIN_XY=6918,8232,6888,8235,6858,8232 $DEVICE_ID=1001
MM512 347 490 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=7707  $PIN_XY=6918,7602,6888,7707,6858,7602 $DEVICE_ID=1001
MM513 GND! 486 98 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6216 $Y=7686  $PIN_XY=6246,7602,6216,7686,6186,7602 $DEVICE_ID=1001
MM514 98 486 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6048 $Y=7686  $PIN_XY=6078,7602,6048,7686,6018,7602 $DEVICE_ID=1001
MM515 GND! 511 486 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5376 $Y=7707  $PIN_XY=5406,7602,5376,7707,5346,7602 $DEVICE_ID=1001
MM516 486 511 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5208 $Y=7707  $PIN_XY=5238,7602,5208,7707,5178,7602 $DEVICE_ID=1001
MM517 GND! 510 469 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5208 $Y=4935  $PIN_XY=5238,4830,5208,4935,5178,4830 $DEVICE_ID=1001
MM518 469 509 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5040 $Y=4914  $PIN_XY=5070,4830,5040,4914,5010,4830 $DEVICE_ID=1001
MM519 485 508 484 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4704 $Y=7707  $PIN_XY=4734,7602,4704,7707,4674,7602 $DEVICE_ID=1001
MM520 484 A<2> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4536 $Y=7707  $PIN_XY=4566,7602,4536,7707,4506,7602 $DEVICE_ID=1001
MM521 GND! 471 96 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4368 $Y=7203  $PIN_XY=4398,7308,4368,7203,4338,7308 $DEVICE_ID=1001
MM522 GND! 469 97 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4368 $Y=4935  $PIN_XY=4398,4830,4368,4935,4338,4830 $DEVICE_ID=1001
MM523 96 471 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4200 $Y=7203  $PIN_XY=4230,7308,4200,7203,4170,7308 $DEVICE_ID=1001
MM524 97 469 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4200 $Y=4935  $PIN_XY=4230,4830,4200,4935,4170,4830 $DEVICE_ID=1001
MM525 83 472 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3696 $Y=4935  $PIN_XY=3726,4830,3696,4935,3666,4830 $DEVICE_ID=1001
MM526 471 507 470 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=7203  $PIN_XY=3390,7308,3360,7203,3330,7308 $DEVICE_ID=1001
MM527 470 506 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=7203  $PIN_XY=3222,7308,3192,7203,3162,7308 $DEVICE_ID=1001
MM528 472 477 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3192 $Y=4914  $PIN_XY=3222,4830,3192,4914,3162,4830 $DEVICE_ID=1001
MM529 477 478 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2688 $Y=4935  $PIN_XY=2718,4830,2688,4935,2658,4830 $DEVICE_ID=1001
MM530 478 475 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2184 $Y=4935  $PIN_XY=2214,4830,2184,4935,2154,4830 $DEVICE_ID=1001
MM531 475 476 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1680 $Y=4935  $PIN_XY=1710,4830,1680,4935,1650,4830 $DEVICE_ID=1001
MM532 476 473 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1176 $Y=4935  $PIN_XY=1206,4830,1176,4935,1146,4830 $DEVICE_ID=1001
MM533 473 474 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=672 $Y=4935  $PIN_XY=702,4830,672,4935,642,4830 $DEVICE_ID=1001
MM534 474 505 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=168 $Y=4935  $PIN_XY=198,4830,168,4935,138,4830 $DEVICE_ID=1001
MM535 94 127 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17472 $Y=1239  $PIN_XY=17502,1134,17472,1239,17442,1134 $DEVICE_ID=1001
MM536 127 24 483 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16968 $Y=1239  $PIN_XY=16998,1134,16968,1239,16938,1134 $DEVICE_ID=1001
MM537 483 338 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16800 $Y=1218  $PIN_XY=16830,1134,16800,1218,16770,1134 $DEVICE_ID=1001
MM538 GND! 73 338 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=1239  $PIN_XY=16158,1134,16128,1239,16098,1134 $DEVICE_ID=1001
MM539 338 73 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=1239  $PIN_XY=15990,1134,15960,1239,15930,1134 $DEVICE_ID=1001
MM540 93 124 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14448 $Y=1239  $PIN_XY=14478,1134,14448,1239,14418,1134 $DEVICE_ID=1001
MM541 124 19 481 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13944 $Y=1239  $PIN_XY=13974,1134,13944,1239,13914,1134 $DEVICE_ID=1001
MM542 481 339 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13776 $Y=1218  $PIN_XY=13806,1134,13776,1218,13746,1134 $DEVICE_ID=1001
MM543 GND! 75 339 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=1239  $PIN_XY=13134,1134,13104,1239,13074,1134 $DEVICE_ID=1001
MM544 339 75 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=1239  $PIN_XY=12966,1134,12936,1239,12906,1134 $DEVICE_ID=1001
MM545 92 121 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11424 $Y=1239  $PIN_XY=11454,1134,11424,1239,11394,1134 $DEVICE_ID=1001
MM546 121 14 482 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10920 $Y=1239  $PIN_XY=10950,1134,10920,1239,10890,1134 $DEVICE_ID=1001
MM547 482 340 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10752 $Y=1218  $PIN_XY=10782,1134,10752,1218,10722,1134 $DEVICE_ID=1001
MM548 GND! 80 340 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=1239  $PIN_XY=10110,1134,10080,1239,10050,1134 $DEVICE_ID=1001
MM549 340 80 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=1239  $PIN_XY=9942,1134,9912,1239,9882,1134 $DEVICE_ID=1001
MM550 91 118 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8400 $Y=1239  $PIN_XY=8430,1134,8400,1239,8370,1134 $DEVICE_ID=1001
MM551 118 9 480 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7896 $Y=1239  $PIN_XY=7926,1134,7896,1239,7866,1134 $DEVICE_ID=1001
MM552 480 328 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7728 $Y=1218  $PIN_XY=7758,1134,7728,1218,7698,1134 $DEVICE_ID=1001
MM553 GND! 78 328 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=1239  $PIN_XY=7086,1134,7056,1239,7026,1134 $DEVICE_ID=1001
MM554 328 78 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=1239  $PIN_XY=6918,1134,6888,1239,6858,1134 $DEVICE_ID=1001
MM555 GND! 89 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6384 $Y=1218  $PIN_XY=6414,1134,6384,1218,6354,1134 $DEVICE_ID=1001
MM556 89 WENB 479 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5880 $Y=1218  $PIN_XY=5910,1134,5880,1218,5850,1134 $DEVICE_ID=1001
MM557 479 83 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5712 $Y=1218  $PIN_XY=5742,1134,5712,1218,5682,1134 $DEVICE_ID=1001
MM558 454 256 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=14154  $PIN_XY=18006,14240,17976,14154,17946,14240 $DEVICE_ID=1003
MM559 452 251 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=13230  $PIN_XY=18006,13316,17976,13230,17946,13316 $DEVICE_ID=1003
MM560 447 245 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=12306  $PIN_XY=18006,12392,17976,12306,17946,12392 $DEVICE_ID=1003
MM561 405 242 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=11382  $PIN_XY=18006,11468,17976,11382,17946,11468 $DEVICE_ID=1003
MM562 402 240 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=10458  $PIN_XY=18006,10544,17976,10458,17946,10544 $DEVICE_ID=1003
MM563 400 170 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=9534  $PIN_XY=18006,9620,17976,9534,17946,9620 $DEVICE_ID=1003
MM564 455 255 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=14154  $PIN_XY=17334,14240,17304,14154,17274,14240 $DEVICE_ID=1003
MM565 451 250 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=13230  $PIN_XY=17334,13316,17304,13230,17274,13316 $DEVICE_ID=1003
MM566 446 246 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=12306  $PIN_XY=17334,12392,17304,12306,17274,12392 $DEVICE_ID=1003
MM567 406 243 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=11382  $PIN_XY=17334,11468,17304,11382,17274,11468 $DEVICE_ID=1003
MM568 403 239 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=10458  $PIN_XY=17334,10544,17304,10458,17274,10544 $DEVICE_ID=1003
MM569 399 172 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=9534  $PIN_XY=17334,9620,17304,9534,17274,9620 $DEVICE_ID=1003
MM570 456 254 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=14154  $PIN_XY=16662,14240,16632,14154,16602,14240 $DEVICE_ID=1003
MM571 450 249 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=13230  $PIN_XY=16662,13316,16632,13230,16602,13316 $DEVICE_ID=1003
MM572 445 247 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=12306  $PIN_XY=16662,12392,16632,12306,16602,12392 $DEVICE_ID=1003
MM573 407 244 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=11382  $PIN_XY=16662,11468,16632,11382,16602,11468 $DEVICE_ID=1003
MM574 404 238 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=10458  $PIN_XY=16662,10544,16632,10458,16602,10544 $DEVICE_ID=1003
MM575 398 174 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=9534  $PIN_XY=16662,9620,16632,9534,16602,9620 $DEVICE_ID=1003
MM576 453 253 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=14154  $PIN_XY=15990,14240,15960,14154,15930,14240 $DEVICE_ID=1003
MM577 449 252 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=13230  $PIN_XY=15990,13316,15960,13230,15930,13316 $DEVICE_ID=1003
MM578 448 248 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=12306  $PIN_XY=15990,12392,15960,12306,15930,12392 $DEVICE_ID=1003
MM579 408 241 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=11382  $PIN_XY=15990,11468,15960,11382,15930,11468 $DEVICE_ID=1003
MM580 401 237 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=10458  $PIN_XY=15990,10544,15960,10458,15930,10544 $DEVICE_ID=1003
MM581 397 176 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=9534  $PIN_XY=15990,9620,15960,9534,15930,9620 $DEVICE_ID=1003
MM582 457 217 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=14154  $PIN_XY=14982,14240,14952,14154,14922,14240 $DEVICE_ID=1003
MM583 458 218 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=13230  $PIN_XY=14982,13316,14952,13230,14922,13316 $DEVICE_ID=1003
MM584 459 219 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=12306  $PIN_XY=14982,12392,14952,12306,14922,12392 $DEVICE_ID=1003
MM585 409 220 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=11382  $PIN_XY=14982,11468,14952,11382,14922,11468 $DEVICE_ID=1003
MM586 410 221 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=10458  $PIN_XY=14982,10544,14952,10458,14922,10544 $DEVICE_ID=1003
MM587 411 158 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=9534  $PIN_XY=14982,9620,14952,9534,14922,9620 $DEVICE_ID=1003
MM588 461 223 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=14154  $PIN_XY=14310,14240,14280,14154,14250,14240 $DEVICE_ID=1003
MM589 463 225 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=13230  $PIN_XY=14310,13316,14280,13230,14250,13316 $DEVICE_ID=1003
MM590 467 229 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=12306  $PIN_XY=14310,12392,14280,12306,14250,12392 $DEVICE_ID=1003
MM591 414 233 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=11382  $PIN_XY=14310,11468,14280,11382,14250,11468 $DEVICE_ID=1003
MM592 416 235 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=10458  $PIN_XY=14310,10544,14280,10458,14250,10544 $DEVICE_ID=1003
MM593 418 164 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=9534  $PIN_XY=14310,9620,14280,9534,14250,9620 $DEVICE_ID=1003
MM594 460 222 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=14154  $PIN_XY=13638,14240,13608,14154,13578,14240 $DEVICE_ID=1003
MM595 464 226 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=13230  $PIN_XY=13638,13316,13608,13230,13578,13316 $DEVICE_ID=1003
MM596 468 230 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=12306  $PIN_XY=13638,12392,13608,12306,13578,12392 $DEVICE_ID=1003
MM597 413 232 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=11382  $PIN_XY=13638,11468,13608,11382,13578,11468 $DEVICE_ID=1003
MM598 415 234 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=10458  $PIN_XY=13638,10544,13608,10458,13578,10544 $DEVICE_ID=1003
MM599 419 162 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=9534  $PIN_XY=13638,9620,13608,9534,13578,9620 $DEVICE_ID=1003
MM600 462 224 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=14154  $PIN_XY=12966,14240,12936,14154,12906,14240 $DEVICE_ID=1003
MM601 465 227 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=13230  $PIN_XY=12966,13316,12936,13230,12906,13316 $DEVICE_ID=1003
MM602 466 228 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=12306  $PIN_XY=12966,12392,12936,12306,12906,12392 $DEVICE_ID=1003
MM603 412 231 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=11382  $PIN_XY=12966,11468,12936,11382,12906,11468 $DEVICE_ID=1003
MM604 417 236 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=10458  $PIN_XY=12966,10544,12936,10458,12906,10544 $DEVICE_ID=1003
MM605 420 160 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=9534  $PIN_XY=12966,9620,12936,9534,12906,9620 $DEVICE_ID=1003
MM606 435 199 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=14154  $PIN_XY=11958,14240,11928,14154,11898,14240 $DEVICE_ID=1003
MM607 437 201 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=13230  $PIN_XY=11958,13316,11928,13230,11898,13316 $DEVICE_ID=1003
MM608 442 206 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=12306  $PIN_XY=11958,12392,11928,12306,11898,12392 $DEVICE_ID=1003
MM609 388 212 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=11382  $PIN_XY=11958,11468,11928,11382,11898,11468 $DEVICE_ID=1003
MM610 391 215 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=10458  $PIN_XY=11958,10544,11928,10458,11898,10544 $DEVICE_ID=1003
MM611 393 152 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=9534  $PIN_XY=11958,9620,11928,9534,11898,9620 $DEVICE_ID=1003
MM612 434 198 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=14154  $PIN_XY=11286,14240,11256,14154,11226,14240 $DEVICE_ID=1003
MM613 438 202 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=13230  $PIN_XY=11286,13316,11256,13230,11226,13316 $DEVICE_ID=1003
MM614 443 207 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=12306  $PIN_XY=11286,12392,11256,12306,11226,12392 $DEVICE_ID=1003
MM615 387 211 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=11382  $PIN_XY=11286,11468,11256,11382,11226,11468 $DEVICE_ID=1003
MM616 390 214 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=10458  $PIN_XY=11286,10544,11256,10458,11226,10544 $DEVICE_ID=1003
MM617 394 150 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=9534  $PIN_XY=11286,9620,11256,9534,11226,9620 $DEVICE_ID=1003
MM618 433 197 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=14154  $PIN_XY=10614,14240,10584,14154,10554,14240 $DEVICE_ID=1003
MM619 439 203 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=13230  $PIN_XY=10614,13316,10584,13230,10554,13316 $DEVICE_ID=1003
MM620 444 208 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=12306  $PIN_XY=10614,12392,10584,12306,10554,12392 $DEVICE_ID=1003
MM621 386 210 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=11382  $PIN_XY=10614,11468,10584,11382,10554,11468 $DEVICE_ID=1003
MM622 389 213 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=10458  $PIN_XY=10614,10544,10584,10458,10554,10544 $DEVICE_ID=1003
MM623 395 148 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=9534  $PIN_XY=10614,9620,10584,9534,10554,9620 $DEVICE_ID=1003
MM624 436 200 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=14154  $PIN_XY=9942,14240,9912,14154,9882,14240 $DEVICE_ID=1003
MM625 440 204 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=13230  $PIN_XY=9942,13316,9912,13230,9882,13316 $DEVICE_ID=1003
MM626 441 205 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=12306  $PIN_XY=9942,12392,9912,12306,9882,12392 $DEVICE_ID=1003
MM627 385 209 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=11382  $PIN_XY=9942,11468,9912,11382,9882,11468 $DEVICE_ID=1003
MM628 392 216 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=10458  $PIN_XY=9942,10544,9912,10458,9882,10544 $DEVICE_ID=1003
MM629 396 146 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=9534  $PIN_XY=9942,9620,9912,9534,9882,9620 $DEVICE_ID=1003
MM630 430 196 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=14154  $PIN_XY=8934,14240,8904,14154,8874,14240 $DEVICE_ID=1003
MM631 428 191 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=13230  $PIN_XY=8934,13316,8904,13230,8874,13316 $DEVICE_ID=1003
MM632 423 185 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=12306  $PIN_XY=8934,12392,8904,12306,8874,12392 $DEVICE_ID=1003
MM633 381 182 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=11382  $PIN_XY=8934,11468,8904,11382,8874,11468 $DEVICE_ID=1003
MM634 378 180 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=10458  $PIN_XY=8934,10544,8904,10458,8874,10544 $DEVICE_ID=1003
MM635 376 138 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=9534  $PIN_XY=8934,9620,8904,9534,8874,9620 $DEVICE_ID=1003
MM636 431 195 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=14154  $PIN_XY=8262,14240,8232,14154,8202,14240 $DEVICE_ID=1003
MM637 427 190 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=13230  $PIN_XY=8262,13316,8232,13230,8202,13316 $DEVICE_ID=1003
MM638 422 186 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=12306  $PIN_XY=8262,12392,8232,12306,8202,12392 $DEVICE_ID=1003
MM639 382 183 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=11382  $PIN_XY=8262,11468,8232,11382,8202,11468 $DEVICE_ID=1003
MM640 379 179 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=10458  $PIN_XY=8262,10544,8232,10458,8202,10544 $DEVICE_ID=1003
MM641 375 137 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=9534  $PIN_XY=8262,9620,8232,9534,8202,9620 $DEVICE_ID=1003
MM642 432 194 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=14154  $PIN_XY=7590,14240,7560,14154,7530,14240 $DEVICE_ID=1003
MM643 426 189 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=13230  $PIN_XY=7590,13316,7560,13230,7530,13316 $DEVICE_ID=1003
MM644 421 187 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=12306  $PIN_XY=7590,12392,7560,12306,7530,12392 $DEVICE_ID=1003
MM645 383 184 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=11382  $PIN_XY=7590,11468,7560,11382,7530,11468 $DEVICE_ID=1003
MM646 380 178 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=10458  $PIN_XY=7590,10544,7560,10458,7530,10544 $DEVICE_ID=1003
MM647 374 136 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=9534  $PIN_XY=7590,9620,7560,9534,7530,9620 $DEVICE_ID=1003
MM648 429 193 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=14154  $PIN_XY=6918,14240,6888,14154,6858,14240 $DEVICE_ID=1003
MM649 425 192 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=13230  $PIN_XY=6918,13316,6888,13230,6858,13316 $DEVICE_ID=1003
MM650 424 188 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=12306  $PIN_XY=6918,12392,6888,12306,6858,12392 $DEVICE_ID=1003
MM651 384 181 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=11382  $PIN_XY=6918,11468,6888,11382,6858,11468 $DEVICE_ID=1003
MM652 377 177 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=10458  $PIN_XY=6918,10544,6888,10458,6858,10544 $DEVICE_ID=1003
MM653 373 140 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=9534  $PIN_XY=6918,9620,6888,9534,6858,9620 $DEVICE_ID=1003
MM654 VDD! 67 27 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18312 $Y=7119  $PIN_XY=18342,7138,18312,7119,18282,7138 $DEVICE_ID=1003
MM655 73 168 27 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18312 $Y=6862  $PIN_XY=18342,6848,18312,6862,18282,6848 $DEVICE_ID=1003
MM656 27 67 24 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18144 $Y=7119  $PIN_XY=18174,7138,18144,7119,18114,7138 $DEVICE_ID=1003
MM657 VDD! WS0 304 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=3528  $PIN_XY=18174,3442,18144,3528,18114,3442 $DEVICE_ID=1003
MM658 357 169 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=8610  $PIN_XY=18006,8696,17976,8610,17946,8696 $DEVICE_ID=1003
MM659 365 500 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=7707  $PIN_XY=18006,7772,17976,7707,17946,7772 $DEVICE_ID=1003
MM660 24 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=7119  $PIN_XY=18006,7138,17976,7119,17946,7138 $DEVICE_ID=1003
MM661 24 168 300 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=6862  $PIN_XY=18006,6848,17976,6862,17946,6848 $DEVICE_ID=1003
MM662 304 82 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=3549  $PIN_XY=18006,3442,17976,3549,17946,3442 $DEVICE_ID=1003
MM663 VDD! 67 26 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17640 $Y=7119  $PIN_XY=17670,7138,17640,7119,17610,7138 $DEVICE_ID=1003
MM664 73 167 26 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17640 $Y=6862  $PIN_XY=17670,6848,17640,6862,17610,6848 $DEVICE_ID=1003
MM665 26 67 24 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17472 $Y=7119  $PIN_XY=17502,7138,17472,7119,17442,7138 $DEVICE_ID=1003
MM666 VDD! 82 303 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=3528  $PIN_XY=17502,3442,17472,3528,17442,3442 $DEVICE_ID=1003
MM667 VDD! 336 72 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=2222  $PIN_XY=17502,2228,17472,2222,17442,2228 $DEVICE_ID=1003
MM668 358 171 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=8610  $PIN_XY=17334,8696,17304,8610,17274,8696 $DEVICE_ID=1003
MM669 364 499 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=7707  $PIN_XY=17334,7772,17304,7707,17274,7772 $DEVICE_ID=1003
MM670 24 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=7119  $PIN_XY=17334,7138,17304,7119,17274,7138 $DEVICE_ID=1003
MM671 24 167 299 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=6862  $PIN_XY=17334,6848,17304,6862,17274,6848 $DEVICE_ID=1003
MM672 303 86 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=3549  $PIN_XY=17334,3442,17304,3549,17274,3442 $DEVICE_ID=1003
MM673 72 336 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17304 $Y=2222  $PIN_XY=17334,2228,17304,2222,17274,2228 $DEVICE_ID=1003
MM674 VDD! 336 72 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17136 $Y=2121  $PIN_XY=17166,2228,17136,2121,17106,2228 $DEVICE_ID=1003
MM675 VDD! 67 25 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16968 $Y=7119  $PIN_XY=16998,7138,16968,7119,16938,7138 $DEVICE_ID=1003
MM676 73 166 25 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16968 $Y=6862  $PIN_XY=16998,6848,16968,6862,16938,6848 $DEVICE_ID=1003
MM677 72 336 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16968 $Y=2121  $PIN_XY=16998,2228,16968,2121,16938,2228 $DEVICE_ID=1003
MM678 25 67 24 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16800 $Y=7119  $PIN_XY=16830,7138,16800,7119,16770,7138 $DEVICE_ID=1003
MM679 VDD! WS0 302 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=3528  $PIN_XY=16830,3442,16800,3528,16770,3442 $DEVICE_ID=1003
MM680 359 173 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=8610  $PIN_XY=16662,8696,16632,8610,16602,8696 $DEVICE_ID=1003
MM681 363 498 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=7707  $PIN_XY=16662,7772,16632,7707,16602,7772 $DEVICE_ID=1003
MM682 24 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=7119  $PIN_XY=16662,7138,16632,7119,16602,7138 $DEVICE_ID=1003
MM683 24 166 73 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=6862  $PIN_XY=16662,6848,16632,6862,16602,6848 $DEVICE_ID=1003
MM684 302 90 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=3549  $PIN_XY=16662,3442,16632,3549,16602,3442 $DEVICE_ID=1003
MM685 VDD! 337 336 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16632 $Y=2222  $PIN_XY=16662,2228,16632,2222,16602,2228 $DEVICE_ID=1003
MM686 336 337 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16464 $Y=2121  $PIN_XY=16494,2228,16464,2121,16434,2228 $DEVICE_ID=1003
MM687 VDD! 67 23 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16296 $Y=7119  $PIN_XY=16326,7138,16296,7119,16266,7138 $DEVICE_ID=1003
MM688 73 165 23 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16296 $Y=6862  $PIN_XY=16326,6848,16296,6862,16266,6848 $DEVICE_ID=1003
MM689 23 67 24 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16128 $Y=7119  $PIN_XY=16158,7138,16128,7119,16098,7138 $DEVICE_ID=1003
MM690 VDD! 90 301 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=3528  $PIN_XY=16158,3442,16128,3528,16098,3442 $DEVICE_ID=1003
MM691 VDD! D<3> 337 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=2222  $PIN_XY=16158,2228,16128,2222,16098,2228 $DEVICE_ID=1003
MM692 360 175 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=8610  $PIN_XY=15990,8696,15960,8610,15930,8696 $DEVICE_ID=1003
MM693 362 497 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=7707  $PIN_XY=15990,7772,15960,7707,15930,7772 $DEVICE_ID=1003
MM694 24 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=7119  $PIN_XY=15990,7138,15960,7119,15930,7138 $DEVICE_ID=1003
MM695 24 165 298 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=6862  $PIN_XY=15990,6848,15960,6862,15930,6848 $DEVICE_ID=1003
MM696 301 86 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=3549  $PIN_XY=15990,3442,15960,3549,15930,3442 $DEVICE_ID=1003
MM697 337 D<3> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=2121  $PIN_XY=15990,2228,15960,2121,15930,2228 $DEVICE_ID=1003
MM698 VDD! 67 22 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15288 $Y=7119  $PIN_XY=15318,7138,15288,7119,15258,7138 $DEVICE_ID=1003
MM699 75 153 22 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15288 $Y=6862  $PIN_XY=15318,6848,15288,6862,15258,6848 $DEVICE_ID=1003
MM700 22 67 19 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=15120 $Y=7119  $PIN_XY=15150,7138,15120,7119,15090,7138 $DEVICE_ID=1003
MM701 VDD! WS0 311 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=3528  $PIN_XY=15150,3442,15120,3528,15090,3442 $DEVICE_ID=1003
MM702 361 157 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=8610  $PIN_XY=14982,8696,14952,8610,14922,8696 $DEVICE_ID=1003
MM703 369 501 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=7707  $PIN_XY=14982,7772,14952,7707,14922,7772 $DEVICE_ID=1003
MM704 19 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=7119  $PIN_XY=14982,7138,14952,7119,14922,7138 $DEVICE_ID=1003
MM705 19 153 307 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=6862  $PIN_XY=14982,6848,14952,6862,14922,6848 $DEVICE_ID=1003
MM706 311 82 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=3549  $PIN_XY=14982,3442,14952,3549,14922,3442 $DEVICE_ID=1003
MM707 VDD! 67 18 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14616 $Y=7119  $PIN_XY=14646,7138,14616,7119,14586,7138 $DEVICE_ID=1003
MM708 75 154 18 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14616 $Y=6862  $PIN_XY=14646,6848,14616,6862,14586,6848 $DEVICE_ID=1003
MM709 18 67 19 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14448 $Y=7119  $PIN_XY=14478,7138,14448,7119,14418,7138 $DEVICE_ID=1003
MM710 VDD! 82 310 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=3528  $PIN_XY=14478,3442,14448,3528,14418,3442 $DEVICE_ID=1003
MM711 VDD! 333 74 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=2222  $PIN_XY=14478,2228,14448,2222,14418,2228 $DEVICE_ID=1003
MM712 368 163 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=8610  $PIN_XY=14310,8696,14280,8610,14250,8696 $DEVICE_ID=1003
MM713 370 502 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=7707  $PIN_XY=14310,7772,14280,7707,14250,7772 $DEVICE_ID=1003
MM714 19 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=7119  $PIN_XY=14310,7138,14280,7119,14250,7138 $DEVICE_ID=1003
MM715 19 154 306 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=6862  $PIN_XY=14310,6848,14280,6862,14250,6848 $DEVICE_ID=1003
MM716 310 86 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=3549  $PIN_XY=14310,3442,14280,3549,14250,3442 $DEVICE_ID=1003
MM717 74 333 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14280 $Y=2222  $PIN_XY=14310,2228,14280,2222,14250,2228 $DEVICE_ID=1003
MM718 VDD! 333 74 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14112 $Y=2121  $PIN_XY=14142,2228,14112,2121,14082,2228 $DEVICE_ID=1003
MM719 VDD! 67 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13944 $Y=7119  $PIN_XY=13974,7138,13944,7119,13914,7138 $DEVICE_ID=1003
MM720 75 155 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13944 $Y=6862  $PIN_XY=13974,6848,13944,6862,13914,6848 $DEVICE_ID=1003
MM721 74 333 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13944 $Y=2121  $PIN_XY=13974,2228,13944,2121,13914,2228 $DEVICE_ID=1003
MM722 20 67 19 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13776 $Y=7119  $PIN_XY=13806,7138,13776,7119,13746,7138 $DEVICE_ID=1003
MM723 VDD! WS0 309 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=3528  $PIN_XY=13806,3442,13776,3528,13746,3442 $DEVICE_ID=1003
MM724 367 161 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=8610  $PIN_XY=13638,8696,13608,8610,13578,8696 $DEVICE_ID=1003
MM725 371 495 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=7707  $PIN_XY=13638,7772,13608,7707,13578,7772 $DEVICE_ID=1003
MM726 19 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=7119  $PIN_XY=13638,7138,13608,7119,13578,7138 $DEVICE_ID=1003
MM727 19 155 75 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=6862  $PIN_XY=13638,6848,13608,6862,13578,6848 $DEVICE_ID=1003
MM728 309 90 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=3549  $PIN_XY=13638,3442,13608,3549,13578,3442 $DEVICE_ID=1003
MM729 VDD! 334 333 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13608 $Y=2222  $PIN_XY=13638,2228,13608,2222,13578,2228 $DEVICE_ID=1003
MM730 333 334 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13440 $Y=2121  $PIN_XY=13470,2228,13440,2121,13410,2228 $DEVICE_ID=1003
MM731 VDD! 67 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13272 $Y=7119  $PIN_XY=13302,7138,13272,7119,13242,7138 $DEVICE_ID=1003
MM732 75 156 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13272 $Y=6862  $PIN_XY=13302,6848,13272,6862,13242,6848 $DEVICE_ID=1003
MM733 21 67 19 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13104 $Y=7119  $PIN_XY=13134,7138,13104,7119,13074,7138 $DEVICE_ID=1003
MM734 VDD! 90 308 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=3528  $PIN_XY=13134,3442,13104,3528,13074,3442 $DEVICE_ID=1003
MM735 VDD! D<2> 334 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=2222  $PIN_XY=13134,2228,13104,2222,13074,2228 $DEVICE_ID=1003
MM736 366 159 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=8610  $PIN_XY=12966,8696,12936,8610,12906,8696 $DEVICE_ID=1003
MM737 372 496 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=7707  $PIN_XY=12966,7772,12936,7707,12906,7772 $DEVICE_ID=1003
MM738 19 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=7119  $PIN_XY=12966,7138,12936,7119,12906,7138 $DEVICE_ID=1003
MM739 19 156 305 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=6862  $PIN_XY=12966,6848,12936,6862,12906,6848 $DEVICE_ID=1003
MM740 308 86 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=3549  $PIN_XY=12966,3442,12936,3549,12906,3442 $DEVICE_ID=1003
MM741 334 D<2> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=2121  $PIN_XY=12966,2228,12936,2121,12906,2228 $DEVICE_ID=1003
MM742 VDD! 67 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12264 $Y=7119  $PIN_XY=12294,7138,12264,7119,12234,7138 $DEVICE_ID=1003
MM743 80 141 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12264 $Y=6862  $PIN_XY=12294,6848,12264,6862,12234,6848 $DEVICE_ID=1003
MM744 17 67 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=12096 $Y=7119  $PIN_XY=12126,7138,12096,7119,12066,7138 $DEVICE_ID=1003
MM745 VDD! WS0 324 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=3528  $PIN_XY=12126,3442,12096,3528,12066,3442 $DEVICE_ID=1003
MM746 352 151 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=8610  $PIN_XY=11958,8696,11928,8610,11898,8696 $DEVICE_ID=1003
MM747 353 491 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=7707  $PIN_XY=11958,7772,11928,7707,11898,7772 $DEVICE_ID=1003
MM748 14 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=7119  $PIN_XY=11958,7138,11928,7119,11898,7138 $DEVICE_ID=1003
MM749 14 141 320 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=6862  $PIN_XY=11958,6848,11928,6862,11898,6848 $DEVICE_ID=1003
MM750 324 82 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=3549  $PIN_XY=11958,3442,11928,3549,11898,3442 $DEVICE_ID=1003
MM751 VDD! 67 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11592 $Y=7119  $PIN_XY=11622,7138,11592,7119,11562,7138 $DEVICE_ID=1003
MM752 80 142 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11592 $Y=6862  $PIN_XY=11622,6848,11592,6862,11562,6848 $DEVICE_ID=1003
MM753 16 67 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11424 $Y=7119  $PIN_XY=11454,7138,11424,7119,11394,7138 $DEVICE_ID=1003
MM754 VDD! 82 323 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=3528  $PIN_XY=11454,3442,11424,3528,11394,3442 $DEVICE_ID=1003
MM755 VDD! 330 79 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=2222  $PIN_XY=11454,2228,11424,2222,11394,2228 $DEVICE_ID=1003
MM756 351 149 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=8610  $PIN_XY=11286,8696,11256,8610,11226,8696 $DEVICE_ID=1003
MM757 354 492 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=7707  $PIN_XY=11286,7772,11256,7707,11226,7772 $DEVICE_ID=1003
MM758 14 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=7119  $PIN_XY=11286,7138,11256,7119,11226,7138 $DEVICE_ID=1003
MM759 14 142 319 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=6862  $PIN_XY=11286,6848,11256,6862,11226,6848 $DEVICE_ID=1003
MM760 323 86 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=3549  $PIN_XY=11286,3442,11256,3549,11226,3442 $DEVICE_ID=1003
MM761 79 330 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11256 $Y=2222  $PIN_XY=11286,2228,11256,2222,11226,2228 $DEVICE_ID=1003
MM762 VDD! 330 79 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11088 $Y=2121  $PIN_XY=11118,2228,11088,2121,11058,2228 $DEVICE_ID=1003
MM763 VDD! 67 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10920 $Y=7119  $PIN_XY=10950,7138,10920,7119,10890,7138 $DEVICE_ID=1003
MM764 80 143 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10920 $Y=6862  $PIN_XY=10950,6848,10920,6862,10890,6848 $DEVICE_ID=1003
MM765 79 330 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10920 $Y=2121  $PIN_XY=10950,2228,10920,2121,10890,2228 $DEVICE_ID=1003
MM766 15 67 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10752 $Y=7119  $PIN_XY=10782,7138,10752,7119,10722,7138 $DEVICE_ID=1003
MM767 VDD! WS0 322 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=3528  $PIN_XY=10782,3442,10752,3528,10722,3442 $DEVICE_ID=1003
MM768 350 147 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=8610  $PIN_XY=10614,8696,10584,8610,10554,8696 $DEVICE_ID=1003
MM769 355 493 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=7707  $PIN_XY=10614,7772,10584,7707,10554,7772 $DEVICE_ID=1003
MM770 14 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=7119  $PIN_XY=10614,7138,10584,7119,10554,7138 $DEVICE_ID=1003
MM771 14 143 80 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=6862  $PIN_XY=10614,6848,10584,6862,10554,6848 $DEVICE_ID=1003
MM772 322 90 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=3549  $PIN_XY=10614,3442,10584,3549,10554,3442 $DEVICE_ID=1003
MM773 VDD! 331 330 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10584 $Y=2222  $PIN_XY=10614,2228,10584,2222,10554,2228 $DEVICE_ID=1003
MM774 330 331 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10416 $Y=2121  $PIN_XY=10446,2228,10416,2121,10386,2228 $DEVICE_ID=1003
MM775 VDD! 67 13 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10248 $Y=7119  $PIN_XY=10278,7138,10248,7119,10218,7138 $DEVICE_ID=1003
MM776 80 144 13 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10248 $Y=6862  $PIN_XY=10278,6848,10248,6862,10218,6848 $DEVICE_ID=1003
MM777 13 67 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10080 $Y=7119  $PIN_XY=10110,7138,10080,7119,10050,7138 $DEVICE_ID=1003
MM778 VDD! 90 321 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=3528  $PIN_XY=10110,3442,10080,3528,10050,3442 $DEVICE_ID=1003
MM779 VDD! D<1> 331 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=2222  $PIN_XY=10110,2228,10080,2222,10050,2228 $DEVICE_ID=1003
MM780 349 145 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=8610  $PIN_XY=9942,8696,9912,8610,9882,8696 $DEVICE_ID=1003
MM781 356 494 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=7707  $PIN_XY=9942,7772,9912,7707,9882,7772 $DEVICE_ID=1003
MM782 14 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=7119  $PIN_XY=9942,7138,9912,7119,9882,7138 $DEVICE_ID=1003
MM783 14 144 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=6862  $PIN_XY=9942,6848,9912,6862,9882,6848 $DEVICE_ID=1003
MM784 321 86 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=3549  $PIN_XY=9942,3442,9912,3549,9882,3442 $DEVICE_ID=1003
MM785 331 D<1> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=2121  $PIN_XY=9942,2228,9912,2121,9882,2228 $DEVICE_ID=1003
MM786 VDD! 67 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9240 $Y=7119  $PIN_XY=9270,7138,9240,7119,9210,7138 $DEVICE_ID=1003
MM787 78 129 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9240 $Y=6862  $PIN_XY=9270,6848,9240,6862,9210,6848 $DEVICE_ID=1003
MM788 8 67 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9072 $Y=7119  $PIN_XY=9102,7138,9072,7119,9042,7138 $DEVICE_ID=1003
MM789 VDD! WS0 318 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=3528  $PIN_XY=9102,3442,9072,3528,9042,3442 $DEVICE_ID=1003
MM790 346 133 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=8610  $PIN_XY=8934,8696,8904,8610,8874,8696 $DEVICE_ID=1003
MM791 341 487 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=7707  $PIN_XY=8934,7772,8904,7707,8874,7772 $DEVICE_ID=1003
MM792 9 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=7119  $PIN_XY=8934,7138,8904,7119,8874,7138 $DEVICE_ID=1003
MM793 9 129 314 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=6862  $PIN_XY=8934,6848,8904,6862,8874,6848 $DEVICE_ID=1003
MM794 318 82 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=3549  $PIN_XY=8934,3442,8904,3549,8874,3442 $DEVICE_ID=1003
MM795 VDD! 67 10 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8568 $Y=7119  $PIN_XY=8598,7138,8568,7119,8538,7138 $DEVICE_ID=1003
MM796 78 130 10 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8568 $Y=6862  $PIN_XY=8598,6848,8568,6862,8538,6848 $DEVICE_ID=1003
MM797 10 67 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8400 $Y=7119  $PIN_XY=8430,7138,8400,7119,8370,7138 $DEVICE_ID=1003
MM798 VDD! 82 317 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=3528  $PIN_XY=8430,3442,8400,3528,8370,3442 $DEVICE_ID=1003
MM799 VDD! 326 77 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=2222  $PIN_XY=8430,2228,8400,2222,8370,2228 $DEVICE_ID=1003
MM800 345 134 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=8610  $PIN_XY=8262,8696,8232,8610,8202,8696 $DEVICE_ID=1003
MM801 342 488 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=7707  $PIN_XY=8262,7772,8232,7707,8202,7772 $DEVICE_ID=1003
MM802 9 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=7119  $PIN_XY=8262,7138,8232,7119,8202,7138 $DEVICE_ID=1003
MM803 9 130 313 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=6862  $PIN_XY=8262,6848,8232,6862,8202,6848 $DEVICE_ID=1003
MM804 317 86 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=3549  $PIN_XY=8262,3442,8232,3549,8202,3442 $DEVICE_ID=1003
MM805 77 326 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8232 $Y=2222  $PIN_XY=8262,2228,8232,2222,8202,2228 $DEVICE_ID=1003
MM806 VDD! 326 77 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8064 $Y=2121  $PIN_XY=8094,2228,8064,2121,8034,2228 $DEVICE_ID=1003
MM807 VDD! 67 11 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7896 $Y=7119  $PIN_XY=7926,7138,7896,7119,7866,7138 $DEVICE_ID=1003
MM808 78 131 11 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7896 $Y=6862  $PIN_XY=7926,6848,7896,6862,7866,6848 $DEVICE_ID=1003
MM809 77 326 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7896 $Y=2121  $PIN_XY=7926,2228,7896,2121,7866,2228 $DEVICE_ID=1003
MM810 11 67 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7728 $Y=7119  $PIN_XY=7758,7138,7728,7119,7698,7138 $DEVICE_ID=1003
MM811 VDD! WS0 316 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=3528  $PIN_XY=7758,3442,7728,3528,7698,3442 $DEVICE_ID=1003
MM812 344 135 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=8610  $PIN_XY=7590,8696,7560,8610,7530,8696 $DEVICE_ID=1003
MM813 343 489 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=7707  $PIN_XY=7590,7772,7560,7707,7530,7772 $DEVICE_ID=1003
MM814 9 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=7119  $PIN_XY=7590,7138,7560,7119,7530,7138 $DEVICE_ID=1003
MM815 9 131 78 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=6862  $PIN_XY=7590,6848,7560,6862,7530,6848 $DEVICE_ID=1003
MM816 316 90 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=3549  $PIN_XY=7590,3442,7560,3549,7530,3442 $DEVICE_ID=1003
MM817 VDD! 327 326 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7560 $Y=2222  $PIN_XY=7590,2228,7560,2222,7530,2228 $DEVICE_ID=1003
MM818 326 327 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7392 $Y=2121  $PIN_XY=7422,2228,7392,2121,7362,2228 $DEVICE_ID=1003
MM819 VDD! 67 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7224 $Y=7119  $PIN_XY=7254,7138,7224,7119,7194,7138 $DEVICE_ID=1003
MM820 78 132 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7224 $Y=6862  $PIN_XY=7254,6848,7224,6862,7194,6848 $DEVICE_ID=1003
MM821 12 67 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7056 $Y=7119  $PIN_XY=7086,7138,7056,7119,7026,7138 $DEVICE_ID=1003
MM822 VDD! 90 315 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=3528  $PIN_XY=7086,3442,7056,3528,7026,3442 $DEVICE_ID=1003
MM823 VDD! D<0> 327 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=2222  $PIN_XY=7086,2228,7056,2222,7026,2228 $DEVICE_ID=1003
MM824 348 139 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=8610  $PIN_XY=6918,8696,6888,8610,6858,8696 $DEVICE_ID=1003
MM825 347 490 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=7707  $PIN_XY=6918,7772,6888,7707,6858,7772 $DEVICE_ID=1003
MM826 9 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=7119  $PIN_XY=6918,7138,6888,7119,6858,7138 $DEVICE_ID=1003
MM827 9 132 312 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=6862  $PIN_XY=6918,6848,6888,6862,6858,6848 $DEVICE_ID=1003
MM828 315 86 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=3549  $PIN_XY=6918,3442,6888,3549,6858,3442 $DEVICE_ID=1003
MM829 327 D<0> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=2121  $PIN_XY=6918,2228,6888,2121,6858,2228 $DEVICE_ID=1003
MM830 VDD! 296 100 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6552 $Y=6842  $PIN_XY=6582,6848,6552,6842,6522,6848 $DEVICE_ID=1003
MM831 VDD! 297 86 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6552 $Y=3528  $PIN_XY=6582,3442,6552,3528,6522,3442 $DEVICE_ID=1003
MM832 100 296 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6384 $Y=6762  $PIN_XY=6414,6848,6384,6762,6354,6848 $DEVICE_ID=1003
MM833 86 297 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6384 $Y=3448  $PIN_XY=6414,3442,6384,3448,6354,3442 $DEVICE_ID=1003
MM834 VDD! 113 297 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6048 $Y=3528  $PIN_XY=6078,3442,6048,3528,6018,3442 $DEVICE_ID=1003
MM835 296 87 295 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5880 $Y=6741  $PIN_XY=5910,6848,5880,6741,5850,6848 $DEVICE_ID=1003
MM836 297 WS0BAR VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5880 $Y=3549  $PIN_XY=5910,3442,5880,3549,5850,3442 $DEVICE_ID=1003
MM837 295 97 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5712 $Y=6762  $PIN_XY=5742,6848,5712,6762,5682,6848 $DEVICE_ID=1003
MM838 VDD! 291 WS0BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5376 $Y=4070  $PIN_XY=5406,4076,5376,4070,5346,4076 $DEVICE_ID=1003
MM839 WS0BAR 291 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5208 $Y=4070  $PIN_XY=5238,4076,5208,4070,5178,4076 $DEVICE_ID=1003
MM840 VDD! 291 WS0BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5040 $Y=3969  $PIN_XY=5070,4076,5040,3969,5010,4076 $DEVICE_ID=1003
MM841 WS0BAR 291 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4872 $Y=3969  $PIN_XY=4902,4076,4872,3969,4842,4076 $DEVICE_ID=1003
MM842 VDD! 503 291 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4368 $Y=3969  $PIN_XY=4398,4076,4368,3969,4338,4076 $DEVICE_ID=1003
MM843 291 288 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4200 $Y=3969  $PIN_XY=4230,4076,4200,3969,4170,4076 $DEVICE_ID=1003
MM844 VDD! 293 288 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=4070  $PIN_XY=3390,4076,3360,4070,3330,4076 $DEVICE_ID=1003
MM845 288 293 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=3990  $PIN_XY=3222,4076,3192,3990,3162,4076 $DEVICE_ID=1003
MM846 VDD! 294 293 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2856 $Y=4070  $PIN_XY=2886,4076,2856,4070,2826,4076 $DEVICE_ID=1003
MM847 293 294 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2688 $Y=3969  $PIN_XY=2718,4076,2688,3969,2658,4076 $DEVICE_ID=1003
MM848 VDD! 292 294 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2184 $Y=3969  $PIN_XY=2214,4076,2184,3969,2154,4076 $DEVICE_ID=1003
MM849 294 A<0> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2016 $Y=3969  $PIN_XY=2046,4076,2016,3969,1986,4076 $DEVICE_ID=1003
MM850 VDD! WENB 292 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1680 $Y=4070  $PIN_XY=1710,4076,1680,4070,1650,4076 $DEVICE_ID=1003
MM851 292 WENB VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1512 $Y=3990  $PIN_XY=1542,4076,1512,3990,1482,4076 $DEVICE_ID=1003
MM852 VDD! 335 66 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18312 $Y=1600  $PIN_XY=18342,1594,18312,1600,18282,1594 $DEVICE_ID=1003
MM853 66 335 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18144 $Y=1600  $PIN_XY=18174,1594,18144,1600,18114,1594 $DEVICE_ID=1003
MM854 VDD! 335 66 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17976 $Y=1680  $PIN_XY=18006,1594,17976,1680,17946,1594 $DEVICE_ID=1003
MM855 66 335 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17808 $Y=1680  $PIN_XY=17838,1594,17808,1680,17778,1594 $DEVICE_ID=1003
MM856 VDD! 127 94 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17640 $Y=1298  $PIN_XY=17670,1304,17640,1298,17610,1304 $DEVICE_ID=1003
MM857 VDD! 128 335 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=1579  $PIN_XY=17502,1594,17472,1579,17442,1594 $DEVICE_ID=1003
MM858 94 127 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17472 $Y=1239  $PIN_XY=17502,1304,17472,1239,17442,1304 $DEVICE_ID=1003
MM859 335 128 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17304 $Y=1600  $PIN_XY=17334,1594,17304,1600,17274,1594 $DEVICE_ID=1003
MM860 VDD! 128 335 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17136 $Y=1701  $PIN_XY=17166,1594,17136,1701,17106,1594 $DEVICE_ID=1003
MM861 335 128 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16968 $Y=1680  $PIN_XY=16998,1594,16968,1680,16938,1594 $DEVICE_ID=1003
MM862 VDD! 24 127 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16968 $Y=1239  $PIN_XY=16998,1304,16968,1239,16938,1304 $DEVICE_ID=1003
MM863 127 338 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16800 $Y=1218  $PIN_XY=16830,1304,16800,1218,16770,1304 $DEVICE_ID=1003
MM864 VDD! 126 128 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16632 $Y=1600  $PIN_XY=16662,1594,16632,1600,16602,1594 $DEVICE_ID=1003
MM865 128 126 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16464 $Y=1680  $PIN_XY=16494,1594,16464,1680,16434,1594 $DEVICE_ID=1003
MM866 VDD! 73 338 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16464 $Y=1319  $PIN_XY=16494,1304,16464,1319,16434,1304 $DEVICE_ID=1003
MM867 338 73 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16296 $Y=1298  $PIN_XY=16326,1304,16296,1298,16266,1304 $DEVICE_ID=1003
MM868 VDD! D<3> 126 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=1579  $PIN_XY=16158,1594,16128,1579,16098,1594 $DEVICE_ID=1003
MM869 VDD! 73 338 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16128 $Y=1239  $PIN_XY=16158,1304,16128,1239,16098,1304 $DEVICE_ID=1003
MM870 126 D<3> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=1680  $PIN_XY=15990,1594,15960,1680,15930,1594 $DEVICE_ID=1003
MM871 338 73 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=1239  $PIN_XY=15990,1304,15960,1239,15930,1304 $DEVICE_ID=1003
MM872 VDD! 332 65 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15288 $Y=1600  $PIN_XY=15318,1594,15288,1600,15258,1594 $DEVICE_ID=1003
MM873 65 332 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=15120 $Y=1600  $PIN_XY=15150,1594,15120,1600,15090,1594 $DEVICE_ID=1003
MM874 VDD! 332 65 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14952 $Y=1680  $PIN_XY=14982,1594,14952,1680,14922,1594 $DEVICE_ID=1003
MM875 65 332 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14784 $Y=1680  $PIN_XY=14814,1594,14784,1680,14754,1594 $DEVICE_ID=1003
MM876 VDD! 124 93 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14616 $Y=1298  $PIN_XY=14646,1304,14616,1298,14586,1304 $DEVICE_ID=1003
MM877 VDD! 125 332 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=1579  $PIN_XY=14478,1594,14448,1579,14418,1594 $DEVICE_ID=1003
MM878 93 124 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14448 $Y=1239  $PIN_XY=14478,1304,14448,1239,14418,1304 $DEVICE_ID=1003
MM879 332 125 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14280 $Y=1600  $PIN_XY=14310,1594,14280,1600,14250,1594 $DEVICE_ID=1003
MM880 VDD! 125 332 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14112 $Y=1701  $PIN_XY=14142,1594,14112,1701,14082,1594 $DEVICE_ID=1003
MM881 332 125 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13944 $Y=1680  $PIN_XY=13974,1594,13944,1680,13914,1594 $DEVICE_ID=1003
MM882 VDD! 19 124 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13944 $Y=1239  $PIN_XY=13974,1304,13944,1239,13914,1304 $DEVICE_ID=1003
MM883 124 339 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13776 $Y=1218  $PIN_XY=13806,1304,13776,1218,13746,1304 $DEVICE_ID=1003
MM884 VDD! 123 125 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13608 $Y=1600  $PIN_XY=13638,1594,13608,1600,13578,1594 $DEVICE_ID=1003
MM885 125 123 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13440 $Y=1680  $PIN_XY=13470,1594,13440,1680,13410,1594 $DEVICE_ID=1003
MM886 VDD! 75 339 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13440 $Y=1319  $PIN_XY=13470,1304,13440,1319,13410,1304 $DEVICE_ID=1003
MM887 339 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13272 $Y=1298  $PIN_XY=13302,1304,13272,1298,13242,1304 $DEVICE_ID=1003
MM888 VDD! D<2> 123 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=1579  $PIN_XY=13134,1594,13104,1579,13074,1594 $DEVICE_ID=1003
MM889 VDD! 75 339 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13104 $Y=1239  $PIN_XY=13134,1304,13104,1239,13074,1304 $DEVICE_ID=1003
MM890 123 D<2> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=1680  $PIN_XY=12966,1594,12936,1680,12906,1594 $DEVICE_ID=1003
MM891 339 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=1239  $PIN_XY=12966,1304,12936,1239,12906,1304 $DEVICE_ID=1003
MM892 VDD! 329 64 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12264 $Y=1600  $PIN_XY=12294,1594,12264,1600,12234,1594 $DEVICE_ID=1003
MM893 64 329 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=12096 $Y=1600  $PIN_XY=12126,1594,12096,1600,12066,1594 $DEVICE_ID=1003
MM894 VDD! 329 64 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11928 $Y=1680  $PIN_XY=11958,1594,11928,1680,11898,1594 $DEVICE_ID=1003
MM895 64 329 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11760 $Y=1680  $PIN_XY=11790,1594,11760,1680,11730,1594 $DEVICE_ID=1003
MM896 VDD! 121 92 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11592 $Y=1298  $PIN_XY=11622,1304,11592,1298,11562,1304 $DEVICE_ID=1003
MM897 VDD! 122 329 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=1579  $PIN_XY=11454,1594,11424,1579,11394,1594 $DEVICE_ID=1003
MM898 92 121 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11424 $Y=1239  $PIN_XY=11454,1304,11424,1239,11394,1304 $DEVICE_ID=1003
MM899 329 122 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11256 $Y=1600  $PIN_XY=11286,1594,11256,1600,11226,1594 $DEVICE_ID=1003
MM900 VDD! 122 329 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11088 $Y=1701  $PIN_XY=11118,1594,11088,1701,11058,1594 $DEVICE_ID=1003
MM901 329 122 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10920 $Y=1680  $PIN_XY=10950,1594,10920,1680,10890,1594 $DEVICE_ID=1003
MM902 VDD! 14 121 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10920 $Y=1239  $PIN_XY=10950,1304,10920,1239,10890,1304 $DEVICE_ID=1003
MM903 121 340 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10752 $Y=1218  $PIN_XY=10782,1304,10752,1218,10722,1304 $DEVICE_ID=1003
MM904 VDD! 120 122 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10584 $Y=1600  $PIN_XY=10614,1594,10584,1600,10554,1594 $DEVICE_ID=1003
MM905 122 120 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10416 $Y=1680  $PIN_XY=10446,1594,10416,1680,10386,1594 $DEVICE_ID=1003
MM906 VDD! 80 340 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10416 $Y=1319  $PIN_XY=10446,1304,10416,1319,10386,1304 $DEVICE_ID=1003
MM907 340 80 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10248 $Y=1298  $PIN_XY=10278,1304,10248,1298,10218,1304 $DEVICE_ID=1003
MM908 VDD! D<1> 120 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=1579  $PIN_XY=10110,1594,10080,1579,10050,1594 $DEVICE_ID=1003
MM909 VDD! 80 340 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10080 $Y=1239  $PIN_XY=10110,1304,10080,1239,10050,1304 $DEVICE_ID=1003
MM910 120 D<1> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=1680  $PIN_XY=9942,1594,9912,1680,9882,1594 $DEVICE_ID=1003
MM911 340 80 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=1239  $PIN_XY=9942,1304,9912,1239,9882,1304 $DEVICE_ID=1003
MM912 VDD! 325 63 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9240 $Y=1600  $PIN_XY=9270,1594,9240,1600,9210,1594 $DEVICE_ID=1003
MM913 63 325 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9072 $Y=1600  $PIN_XY=9102,1594,9072,1600,9042,1594 $DEVICE_ID=1003
MM914 VDD! 325 63 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8904 $Y=1680  $PIN_XY=8934,1594,8904,1680,8874,1594 $DEVICE_ID=1003
MM915 63 325 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8736 $Y=1680  $PIN_XY=8766,1594,8736,1680,8706,1594 $DEVICE_ID=1003
MM916 VDD! 118 91 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8568 $Y=1298  $PIN_XY=8598,1304,8568,1298,8538,1304 $DEVICE_ID=1003
MM917 VDD! 119 325 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=1579  $PIN_XY=8430,1594,8400,1579,8370,1594 $DEVICE_ID=1003
MM918 91 118 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8400 $Y=1239  $PIN_XY=8430,1304,8400,1239,8370,1304 $DEVICE_ID=1003
MM919 325 119 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8232 $Y=1600  $PIN_XY=8262,1594,8232,1600,8202,1594 $DEVICE_ID=1003
MM920 VDD! 119 325 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8064 $Y=1701  $PIN_XY=8094,1594,8064,1701,8034,1594 $DEVICE_ID=1003
MM921 325 119 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7896 $Y=1680  $PIN_XY=7926,1594,7896,1680,7866,1594 $DEVICE_ID=1003
MM922 VDD! 9 118 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7896 $Y=1239  $PIN_XY=7926,1304,7896,1239,7866,1304 $DEVICE_ID=1003
MM923 118 328 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7728 $Y=1218  $PIN_XY=7758,1304,7728,1218,7698,1304 $DEVICE_ID=1003
MM924 VDD! 117 119 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7560 $Y=1600  $PIN_XY=7590,1594,7560,1600,7530,1594 $DEVICE_ID=1003
MM925 119 117 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7392 $Y=1680  $PIN_XY=7422,1594,7392,1680,7362,1594 $DEVICE_ID=1003
MM926 VDD! 78 328 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7392 $Y=1319  $PIN_XY=7422,1304,7392,1319,7362,1304 $DEVICE_ID=1003
MM927 328 78 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7224 $Y=1298  $PIN_XY=7254,1304,7224,1298,7194,1304 $DEVICE_ID=1003
MM928 VDD! D<0> 117 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=1579  $PIN_XY=7086,1594,7056,1579,7026,1594 $DEVICE_ID=1003
MM929 VDD! 78 328 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7056 $Y=1239  $PIN_XY=7086,1304,7056,1239,7026,1304 $DEVICE_ID=1003
MM930 117 D<0> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=1680  $PIN_XY=6918,1594,6888,1680,6858,1594 $DEVICE_ID=1003
MM931 328 78 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=1239  $PIN_XY=6918,1304,6888,1239,6858,1304 $DEVICE_ID=1003
MM932 VDD! 89 GND! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6552 $Y=1298  $PIN_XY=6582,1304,6552,1298,6522,1304 $DEVICE_ID=1003
MM933 GND! 89 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6384 $Y=1218  $PIN_XY=6414,1304,6384,1218,6354,1304 $DEVICE_ID=1003
MM934 VDD! WENB 89 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5880 $Y=1218  $PIN_XY=5910,1304,5880,1218,5850,1304 $DEVICE_ID=1003
MM935 89 83 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5712 $Y=1218  $PIN_XY=5742,1304,5712,1218,5682,1304 $DEVICE_ID=1003
MM936 VDD! 290 70 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5376 $Y=676  $PIN_XY=5406,670,5376,676,5346,670 $DEVICE_ID=1003
MM937 70 290 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5208 $Y=676  $PIN_XY=5238,670,5208,676,5178,670 $DEVICE_ID=1003
MM938 VDD! 290 70 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5040 $Y=777  $PIN_XY=5070,670,5040,777,5010,670 $DEVICE_ID=1003
MM939 70 290 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4872 $Y=777  $PIN_XY=4902,670,4872,777,4842,670 $DEVICE_ID=1003
MM940 VDD! 504 289 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4536 $Y=777  $PIN_XY=4566,670,4536,777,4506,670 $DEVICE_ID=1003
MM941 289 503 290 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4368 $Y=777  $PIN_XY=4398,670,4368,777,4338,670 $DEVICE_ID=1003
XX30BB92C51 GND! VDD! GND! 89 257 277 inv $T=6162 924 0 0 $X=6162 $Y=924
XX30BB92C52 VDD! GND! VDD! D<0> 119 326 77 63 117 327 78 
+	78 78 118 _GENERATED_544 _GENERATED_546 _GENERATED_545 _GENERATED_547 9 259 277 278 
+	325 Write_Driver $T=6518 828 0 0 $X=6665 $Y=1384
XX30BB92C53 VDD! GND! VDD! D<1> 122 330 79 64 120 331 80 
+	80 80 121 _GENERATED_548 _GENERATED_550 _GENERATED_549 _GENERATED_551 14 259 277 278 
+	329 Write_Driver $T=9542 828 0 0 $X=9690 $Y=1384
XX30BB92C54 VDD! GND! VDD! D<2> 125 333 74 65 123 334 75 
+	75 75 124 _GENERATED_552 _GENERATED_554 _GENERATED_553 _GENERATED_555 19 259 277 278 
+	332 Write_Driver $T=12566 828 0 0 $X=12714 $Y=1384
XX30BB92C55 VDD! GND! VDD! D<3> 128 336 72 66 126 337 73 
+	73 73 127 VDD! GND! VDD! GND! 24 259 277 278 
+	335 Write_Driver $T=15590 828 0 0 $X=15738 $Y=1384
XX30BB92C56 VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! 293 504 
+	288 WENB 503 291 WS0 70 69 WS1 WS1BAR 87 71 
+	WS0BAR 290 A<1> A<0> 257 258 259 260 277 278 276 
+	275 274 289 292 294 agen_unit $T=1288 2074 0 0 $X=1290 $Y=459
XX30BB92C57 VDD! GND! 8 9 67 129 129 262 VDD! precharge_logic $T=9462 7518 0 180 $X=8682 $Y=6930
XX30BB92C58 VDD! GND! 10 9 67 130 130 262 VDD! precharge_logic $T=8790 7518 0 180 $X=8010 $Y=6930
XX30BB92C59 VDD! GND! 11 9 67 131 131 262 VDD! precharge_logic $T=8118 7518 0 180 $X=7338 $Y=6930
XX30BB92C510 VDD! GND! 12 9 67 132 132 262 VDD! precharge_logic $T=7446 7518 0 180 $X=6665 $Y=6930
XX30BB92C511 VDD! GND! 17 14 67 141 141 262 VDD! precharge_logic $T=12486 7518 0 180 $X=11706 $Y=6930
XX30BB92C512 VDD! GND! 16 14 67 142 142 262 VDD! precharge_logic $T=11814 7518 0 180 $X=11034 $Y=6930
XX30BB92C513 VDD! GND! 15 14 67 143 143 262 VDD! precharge_logic $T=11142 7518 0 180 $X=10362 $Y=6930
XX30BB92C514 VDD! GND! 13 14 67 144 144 262 VDD! precharge_logic $T=10470 7518 0 180 $X=9690 $Y=6930
XX30BB92C515 VDD! GND! 23 24 67 165 165 262 VDD! precharge_logic $T=16518 7518 0 180 $X=15738 $Y=6930
XX30BB92C516 VDD! GND! 25 24 67 166 166 262 VDD! precharge_logic $T=17190 7518 0 180 $X=16410 $Y=6930
XX30BB92C517 VDD! GND! 26 24 67 167 167 262 VDD! precharge_logic $T=17862 7518 0 180 $X=17082 $Y=6930
XX30BB92C518 VDD! GND! 27 24 67 168 168 262 VDD! precharge_logic $T=18534 7518 0 180 $X=17753 $Y=6930
XX30BB92C519 VDD! GND! 22 19 67 153 153 262 VDD! precharge_logic $T=15510 7518 0 180 $X=14730 $Y=6930
XX30BB92C520 VDD! GND! 18 19 67 154 154 262 VDD! precharge_logic $T=14838 7518 0 180 $X=14058 $Y=6930
XX30BB92C521 VDD! GND! 20 19 67 155 155 262 VDD! precharge_logic $T=14166 7518 0 180 $X=13386 $Y=6930
XX30BB92C522 VDD! GND! 21 19 67 156 156 262 VDD! precharge_logic $T=13494 7518 0 180 $X=12714 $Y=6930
XX30BB92C523 GND! VDD! 89 83 WENB 479 257 277 nand $T=5072 696 0 0 $X=5490 $Y=924
XX30BB92C524 GND! VDD! VDD! GND! VDD! GND! VDD! GND! VDD! 296 297 
+	97 113 69 70 87 71 WS0BAR WS1 WS0 68 85 
+	86 82 WS1BAR 90 76 100 260 261 263 264 275 
+	274 279 VDD! VDD! 295 between_blocks $T=5162 4502 0 0 $X=5490 $Y=3231
XX30BB92C525 GND! VDD! GND! VDD! VDD! GND! GND! 505 473 506 475 
+	507 510 CLK 477 471 83 469 509 96 97 67 
+	472 474 476 478 262 264 263 261 VDD! 279 VDD! 
+	470 WLRef_PC $T=-394 4618 0 0 $X=-53 $Y=4620
XX30BB92C526 GND! VDD! _GENERATED_557 _GENERATED_556 47 48 271 285 Filler $T=-58 14910 1 0 $X=-54 $Y=14320
XX30BB92C527 GND! VDD! _GENERATED_559 _GENERATED_558 49 50 270 285 Filler $T=-58 13860 0 0 $X=-54 $Y=13860
XX30BB92C528 GND! VDD! _GENERATED_561 _GENERATED_560 51 52 270 286 Filler $T=-58 13986 1 0 $X=-54 $Y=13396
XX30BB92C529 GND! VDD! _GENERATED_563 _GENERATED_562 53 54 269 286 Filler $T=-58 12936 0 0 $X=-54 $Y=12936
XX30BB92C530 GND! VDD! _GENERATED_565 _GENERATED_564 55 56 268 287 Filler $T=-58 12012 0 0 $X=-54 $Y=12012
XX30BB92C531 GND! VDD! _GENERATED_567 _GENERATED_566 57 58 269 287 Filler $T=-58 13062 1 0 $X=-54 $Y=12472
XX30BB92C532 GND! VDD! _GENERATED_569 _GENERATED_568 31 32 267 283 Filler $T=-58 11088 0 0 $X=-54 $Y=11088
XX30BB92C533 GND! VDD! _GENERATED_571 _GENERATED_570 59 60 268 283 Filler $T=-58 12138 1 0 $X=-54 $Y=11548
XX30BB92C534 GND! VDD! _GENERATED_573 _GENERATED_572 33 34 267 284 Filler $T=-58 11214 1 0 $X=-54 $Y=10624
XX30BB92C535 GND! VDD! _GENERATED_575 _GENERATED_574 35 36 266 284 Filler $T=-58 10164 0 0 $X=-54 $Y=10164
XX30BB92C536 GND! VDD! _GENERATED_577 _GENERATED_576 37 38 266 282 Filler $T=-58 10290 1 0 $X=-54 $Y=9700
XX30BB92C537 GND! VDD! _GENERATED_579 _GENERATED_578 39 40 265 282 Filler $T=-58 9240 0 0 $X=-54 $Y=9240
XX30BB92C538 GND! VDD! _GENERATED_581 _GENERATED_580 41 42 265 280 Filler $T=-58 9366 1 0 $X=-54 $Y=8776
XX30BB92C539 GND! VDD! _GENERATED_583 _GENERATED_582 43 44 272 280 Filler $T=-58 8316 0 0 $X=-54 $Y=8316
XX30BB92C540 GND! VDD! _GENERATED_585 _GENERATED_584 45 46 272 281 Filler $T=-58 8442 1 0 $X=-54 $Y=7852
XX30BB92C541 GND! VDD! _GENERATED_587 _GENERATED_586 29 30 262 281 Filler $T=-58 7392 0 0 $X=-54 $Y=7392
XX30BB92C542 GND! VDD! 47 48 _GENERATED_589 _GENERATED_588 271 285 Filler $T=110 14910 1 0 $X=114 $Y=14320
XX30BB92C543 GND! VDD! 49 50 _GENERATED_591 _GENERATED_590 270 285 Filler $T=110 13860 0 0 $X=114 $Y=13860
XX30BB92C544 GND! VDD! 51 52 _GENERATED_593 _GENERATED_592 270 286 Filler $T=110 13986 1 0 $X=114 $Y=13396
XX30BB92C545 GND! VDD! 53 54 _GENERATED_595 _GENERATED_594 269 286 Filler $T=110 12936 0 0 $X=114 $Y=12936
XX30BB92C546 GND! VDD! 55 56 _GENERATED_597 _GENERATED_596 268 287 Filler $T=110 12012 0 0 $X=114 $Y=12012
XX30BB92C547 GND! VDD! 57 58 _GENERATED_599 _GENERATED_598 269 287 Filler $T=110 13062 1 0 $X=114 $Y=12472
XX30BB92C548 GND! VDD! 31 32 _GENERATED_601 _GENERATED_600 267 283 Filler $T=110 11088 0 0 $X=114 $Y=11088
XX30BB92C549 GND! VDD! 59 60 _GENERATED_603 _GENERATED_602 268 283 Filler $T=110 12138 1 0 $X=114 $Y=11548
XX30BB92C550 GND! VDD! 43 44 _GENERATED_605 _GENERATED_604 272 280 Filler $T=110 8316 0 0 $X=114 $Y=8316
XX30BB92C551 GND! VDD! 29 30 _GENERATED_607 _GENERATED_606 262 281 Filler $T=110 7392 0 0 $X=114 $Y=7392
XX30BB92C552 GND! VDD! 45 46 _GENERATED_609 _GENERATED_608 272 281 Filler $T=110 8442 1 0 $X=114 $Y=7852
XX30BB92C553 GND! VDD! 41 42 _GENERATED_611 _GENERATED_610 265 280 Filler $T=110 9366 1 0 $X=114 $Y=8776
XX30BB92C554 GND! VDD! 33 34 _GENERATED_613 _GENERATED_612 267 284 Filler $T=110 11214 1 0 $X=114 $Y=10624
XX30BB92C555 GND! VDD! 35 36 _GENERATED_615 _GENERATED_614 266 284 Filler $T=110 10164 0 0 $X=114 $Y=10164
XX30BB92C556 GND! VDD! 37 38 _GENERATED_617 _GENERATED_616 266 282 Filler $T=110 10290 1 0 $X=114 $Y=9700
XX30BB92C557 GND! VDD! 39 40 _GENERATED_619 _GENERATED_618 265 282 Filler $T=110 9240 0 0 $X=114 $Y=9240
XX30BB92C558 GND! VDD! _GENERATED_622 _GENERATED_620 _GENERATED_623 _GENERATED_621 262 281 Filler $T=446 7392 0 0 $X=450 $Y=7392
XX30BB92C559 GND! VDD! _GENERATED_626 _GENERATED_624 _GENERATED_627 _GENERATED_625 272 281 Filler $T=446 8442 1 0 $X=450 $Y=7852
XX30BB92C560 GND! VDD! _GENERATED_630 _GENERATED_628 _GENERATED_631 _GENERATED_629 272 280 Filler $T=446 8316 0 0 $X=450 $Y=8316
XX30BB92C561 GND! VDD! _GENERATED_634 _GENERATED_632 _GENERATED_635 _GENERATED_633 265 280 Filler $T=446 9366 1 0 $X=450 $Y=8776
XX30BB92C562 GND! VDD! _GENERATED_638 _GENERATED_636 _GENERATED_639 _GENERATED_637 265 282 Filler $T=446 9240 0 0 $X=450 $Y=9240
XX30BB92C563 GND! VDD! _GENERATED_642 _GENERATED_640 _GENERATED_643 _GENERATED_641 266 282 Filler $T=446 10290 1 0 $X=450 $Y=9700
XX30BB92C564 GND! VDD! _GENERATED_646 _GENERATED_644 _GENERATED_647 _GENERATED_645 266 284 Filler $T=446 10164 0 0 $X=450 $Y=10164
XX30BB92C565 GND! VDD! _GENERATED_650 _GENERATED_648 _GENERATED_651 _GENERATED_649 267 284 Filler $T=446 11214 1 0 $X=450 $Y=10624
XX30BB92C566 GND! VDD! _GENERATED_654 _GENERATED_652 _GENERATED_655 _GENERATED_653 268 283 Filler $T=446 12138 1 0 $X=450 $Y=11548
XX30BB92C567 GND! VDD! _GENERATED_658 _GENERATED_656 _GENERATED_659 _GENERATED_657 267 283 Filler $T=446 11088 0 0 $X=450 $Y=11088
XX30BB92C568 GND! VDD! _GENERATED_662 _GENERATED_660 _GENERATED_663 _GENERATED_661 269 287 Filler $T=446 13062 1 0 $X=450 $Y=12472
XX30BB92C569 GND! VDD! _GENERATED_666 _GENERATED_664 _GENERATED_667 _GENERATED_665 268 287 Filler $T=446 12012 0 0 $X=450 $Y=12012
XX30BB92C570 GND! VDD! _GENERATED_670 _GENERATED_668 _GENERATED_671 _GENERATED_669 269 286 Filler $T=446 12936 0 0 $X=450 $Y=12936
XX30BB92C571 GND! VDD! _GENERATED_674 _GENERATED_672 _GENERATED_675 _GENERATED_673 270 286 Filler $T=446 13986 1 0 $X=450 $Y=13396
XX30BB92C572 GND! VDD! _GENERATED_678 _GENERATED_676 _GENERATED_679 _GENERATED_677 270 285 Filler $T=446 13860 0 0 $X=450 $Y=13860
XX30BB92C573 GND! VDD! _GENERATED_682 _GENERATED_680 _GENERATED_683 _GENERATED_681 271 285 Filler $T=446 14910 1 0 $X=450 $Y=14320
XX30BB92C574 GND! VDD! _GENERATED_686 _GENERATED_684 _GENERATED_687 _GENERATED_685 265 282 Filler $T=782 9240 0 0 $X=786 $Y=9240
XX30BB92C575 GND! VDD! _GENERATED_690 _GENERATED_688 _GENERATED_691 _GENERATED_689 266 282 Filler $T=782 10290 1 0 $X=786 $Y=9700
XX30BB92C576 GND! VDD! _GENERATED_694 _GENERATED_692 _GENERATED_695 _GENERATED_693 266 284 Filler $T=782 10164 0 0 $X=786 $Y=10164
XX30BB92C577 GND! VDD! _GENERATED_698 _GENERATED_696 _GENERATED_699 _GENERATED_697 267 284 Filler $T=782 11214 1 0 $X=786 $Y=10624
XX30BB92C578 GND! VDD! _GENERATED_702 _GENERATED_700 _GENERATED_703 _GENERATED_701 265 280 Filler $T=782 9366 1 0 $X=786 $Y=8776
XX30BB92C579 GND! VDD! _GENERATED_706 _GENERATED_704 _GENERATED_707 _GENERATED_705 272 281 Filler $T=782 8442 1 0 $X=786 $Y=7852
XX30BB92C580 GND! VDD! _GENERATED_710 _GENERATED_708 _GENERATED_711 _GENERATED_709 262 281 Filler $T=782 7392 0 0 $X=786 $Y=7392
XX30BB92C581 GND! VDD! _GENERATED_714 _GENERATED_712 _GENERATED_715 _GENERATED_713 272 280 Filler $T=782 8316 0 0 $X=786 $Y=8316
XX30BB92C582 GND! VDD! _GENERATED_718 _GENERATED_716 _GENERATED_719 _GENERATED_717 268 283 Filler $T=782 12138 1 0 $X=786 $Y=11548
XX30BB92C583 GND! VDD! _GENERATED_722 _GENERATED_720 _GENERATED_723 _GENERATED_721 267 283 Filler $T=782 11088 0 0 $X=786 $Y=11088
XX30BB92C584 GND! VDD! _GENERATED_726 _GENERATED_724 _GENERATED_727 _GENERATED_725 269 287 Filler $T=782 13062 1 0 $X=786 $Y=12472
XX30BB92C585 GND! VDD! _GENERATED_730 _GENERATED_728 _GENERATED_731 _GENERATED_729 268 287 Filler $T=782 12012 0 0 $X=786 $Y=12012
XX30BB92C586 GND! VDD! _GENERATED_734 _GENERATED_732 _GENERATED_735 _GENERATED_733 269 286 Filler $T=782 12936 0 0 $X=786 $Y=12936
XX30BB92C587 GND! VDD! _GENERATED_738 _GENERATED_736 _GENERATED_739 _GENERATED_737 270 286 Filler $T=782 13986 1 0 $X=786 $Y=13396
XX30BB92C588 GND! VDD! _GENERATED_742 _GENERATED_740 _GENERATED_743 _GENERATED_741 270 285 Filler $T=782 13860 0 0 $X=786 $Y=13860
XX30BB92C589 GND! VDD! _GENERATED_746 _GENERATED_744 _GENERATED_747 _GENERATED_745 271 285 Filler $T=782 14910 1 0 $X=786 $Y=14320
XX30BB92C590 GND! VDD! _GENERATED_750 _GENERATED_748 _GENERATED_751 _GENERATED_749 271 285 Filler $T=1118 14910 1 0 $X=1122 $Y=14320
XX30BB92C591 GND! VDD! _GENERATED_754 _GENERATED_752 _GENERATED_755 _GENERATED_753 270 285 Filler $T=1118 13860 0 0 $X=1122 $Y=13860
XX30BB92C592 GND! VDD! _GENERATED_758 _GENERATED_756 _GENERATED_759 _GENERATED_757 270 286 Filler $T=1118 13986 1 0 $X=1122 $Y=13396
XX30BB92C593 GND! VDD! _GENERATED_762 _GENERATED_760 _GENERATED_763 _GENERATED_761 269 286 Filler $T=1118 12936 0 0 $X=1122 $Y=12936
XX30BB92C594 GND! VDD! _GENERATED_766 _GENERATED_764 _GENERATED_767 _GENERATED_765 268 287 Filler $T=1118 12012 0 0 $X=1122 $Y=12012
XX30BB92C595 GND! VDD! _GENERATED_770 _GENERATED_768 _GENERATED_771 _GENERATED_769 269 287 Filler $T=1118 13062 1 0 $X=1122 $Y=12472
XX30BB92C596 GND! VDD! _GENERATED_774 _GENERATED_772 _GENERATED_775 _GENERATED_773 267 283 Filler $T=1118 11088 0 0 $X=1122 $Y=11088
XX30BB92C597 GND! VDD! _GENERATED_778 _GENERATED_776 _GENERATED_779 _GENERATED_777 268 283 Filler $T=1118 12138 1 0 $X=1122 $Y=11548
XX30BB92C598 GND! VDD! _GENERATED_782 _GENERATED_780 _GENERATED_783 _GENERATED_781 267 284 Filler $T=1118 11214 1 0 $X=1122 $Y=10624
XX30BB92C599 GND! VDD! _GENERATED_786 _GENERATED_784 _GENERATED_787 _GENERATED_785 266 284 Filler $T=1118 10164 0 0 $X=1122 $Y=10164
XX30BB92C5100 GND! VDD! _GENERATED_790 _GENERATED_788 _GENERATED_791 _GENERATED_789 266 282 Filler $T=1118 10290 1 0 $X=1122 $Y=9700
XX30BB92C5101 GND! VDD! _GENERATED_794 _GENERATED_792 _GENERATED_795 _GENERATED_793 265 282 Filler $T=1118 9240 0 0 $X=1122 $Y=9240
XX30BB92C5102 GND! VDD! _GENERATED_798 _GENERATED_796 _GENERATED_799 _GENERATED_797 265 280 Filler $T=1118 9366 1 0 $X=1122 $Y=8776
XX30BB92C5103 GND! VDD! _GENERATED_802 _GENERATED_800 _GENERATED_803 _GENERATED_801 272 280 Filler $T=1118 8316 0 0 $X=1122 $Y=8316
XX30BB92C5104 GND! VDD! _GENERATED_806 _GENERATED_804 _GENERATED_807 _GENERATED_805 272 281 Filler $T=1118 8442 1 0 $X=1122 $Y=7852
XX30BB92C5105 GND! VDD! _GENERATED_810 _GENERATED_808 _GENERATED_811 _GENERATED_809 262 281 Filler $T=1118 7392 0 0 $X=1122 $Y=7392
XX30BB92C5106 GND! VDD! _GENERATED_814 _GENERATED_812 _GENERATED_815 _GENERATED_813 271 285 Filler $T=1454 14910 1 0 $X=1458 $Y=14320
XX30BB92C5107 GND! VDD! _GENERATED_818 _GENERATED_816 _GENERATED_819 _GENERATED_817 270 285 Filler $T=1454 13860 0 0 $X=1458 $Y=13860
XX30BB92C5108 GND! VDD! _GENERATED_822 _GENERATED_820 _GENERATED_823 _GENERATED_821 270 286 Filler $T=1454 13986 1 0 $X=1458 $Y=13396
XX30BB92C5109 GND! VDD! _GENERATED_826 _GENERATED_824 _GENERATED_827 _GENERATED_825 269 286 Filler $T=1454 12936 0 0 $X=1458 $Y=12936
XX30BB92C5110 GND! VDD! _GENERATED_830 _GENERATED_828 _GENERATED_831 _GENERATED_829 268 287 Filler $T=1454 12012 0 0 $X=1458 $Y=12012
XX30BB92C5111 GND! VDD! _GENERATED_834 _GENERATED_832 _GENERATED_835 _GENERATED_833 269 287 Filler $T=1454 13062 1 0 $X=1458 $Y=12472
XX30BB92C5112 GND! VDD! _GENERATED_838 _GENERATED_836 _GENERATED_839 _GENERATED_837 267 283 Filler $T=1454 11088 0 0 $X=1458 $Y=11088
XX30BB92C5113 GND! VDD! _GENERATED_842 _GENERATED_840 _GENERATED_843 _GENERATED_841 268 283 Filler $T=1454 12138 1 0 $X=1458 $Y=11548
XX30BB92C5114 GND! VDD! _GENERATED_846 _GENERATED_844 _GENERATED_847 _GENERATED_845 272 280 Filler $T=1454 8316 0 0 $X=1458 $Y=8316
XX30BB92C5115 GND! VDD! _GENERATED_850 _GENERATED_848 _GENERATED_851 _GENERATED_849 262 281 Filler $T=1454 7392 0 0 $X=1458 $Y=7392
XX30BB92C5116 GND! VDD! _GENERATED_854 _GENERATED_852 _GENERATED_855 _GENERATED_853 272 281 Filler $T=1454 8442 1 0 $X=1458 $Y=7852
XX30BB92C5117 GND! VDD! _GENERATED_858 _GENERATED_856 _GENERATED_859 _GENERATED_857 265 280 Filler $T=1454 9366 1 0 $X=1458 $Y=8776
XX30BB92C5118 GND! VDD! _GENERATED_862 _GENERATED_860 _GENERATED_863 _GENERATED_861 267 284 Filler $T=1454 11214 1 0 $X=1458 $Y=10624
XX30BB92C5119 GND! VDD! _GENERATED_866 _GENERATED_864 _GENERATED_867 _GENERATED_865 266 284 Filler $T=1454 10164 0 0 $X=1458 $Y=10164
XX30BB92C5120 GND! VDD! _GENERATED_870 _GENERATED_868 _GENERATED_871 _GENERATED_869 266 282 Filler $T=1454 10290 1 0 $X=1458 $Y=9700
XX30BB92C5121 GND! VDD! _GENERATED_874 _GENERATED_872 _GENERATED_875 _GENERATED_873 265 282 Filler $T=1454 9240 0 0 $X=1458 $Y=9240
XX30BB92C5122 GND! VDD! _GENERATED_878 _GENERATED_876 _GENERATED_879 _GENERATED_877 262 281 Filler $T=1790 7392 0 0 $X=1794 $Y=7392
XX30BB92C5123 GND! VDD! _GENERATED_882 _GENERATED_880 _GENERATED_883 _GENERATED_881 272 281 Filler $T=1790 8442 1 0 $X=1794 $Y=7852
XX30BB92C5124 GND! VDD! _GENERATED_886 _GENERATED_884 _GENERATED_887 _GENERATED_885 272 280 Filler $T=1790 8316 0 0 $X=1794 $Y=8316
XX30BB92C5125 GND! VDD! _GENERATED_890 _GENERATED_888 _GENERATED_891 _GENERATED_889 265 280 Filler $T=1790 9366 1 0 $X=1794 $Y=8776
XX30BB92C5126 GND! VDD! _GENERATED_894 _GENERATED_892 _GENERATED_895 _GENERATED_893 265 282 Filler $T=1790 9240 0 0 $X=1794 $Y=9240
XX30BB92C5127 GND! VDD! _GENERATED_898 _GENERATED_896 _GENERATED_899 _GENERATED_897 266 282 Filler $T=1790 10290 1 0 $X=1794 $Y=9700
XX30BB92C5128 GND! VDD! _GENERATED_902 _GENERATED_900 _GENERATED_903 _GENERATED_901 266 284 Filler $T=1790 10164 0 0 $X=1794 $Y=10164
XX30BB92C5129 GND! VDD! _GENERATED_906 _GENERATED_904 _GENERATED_907 _GENERATED_905 267 284 Filler $T=1790 11214 1 0 $X=1794 $Y=10624
XX30BB92C5130 GND! VDD! _GENERATED_910 _GENERATED_908 _GENERATED_911 _GENERATED_909 268 283 Filler $T=1790 12138 1 0 $X=1794 $Y=11548
XX30BB92C5131 GND! VDD! _GENERATED_914 _GENERATED_912 _GENERATED_915 _GENERATED_913 267 283 Filler $T=1790 11088 0 0 $X=1794 $Y=11088
XX30BB92C5132 GND! VDD! _GENERATED_918 _GENERATED_916 _GENERATED_919 _GENERATED_917 269 287 Filler $T=1790 13062 1 0 $X=1794 $Y=12472
XX30BB92C5133 GND! VDD! _GENERATED_922 _GENERATED_920 _GENERATED_923 _GENERATED_921 268 287 Filler $T=1790 12012 0 0 $X=1794 $Y=12012
XX30BB92C5134 GND! VDD! _GENERATED_926 _GENERATED_924 _GENERATED_927 _GENERATED_925 269 286 Filler $T=1790 12936 0 0 $X=1794 $Y=12936
XX30BB92C5135 GND! VDD! _GENERATED_930 _GENERATED_928 _GENERATED_931 _GENERATED_929 270 286 Filler $T=1790 13986 1 0 $X=1794 $Y=13396
XX30BB92C5136 GND! VDD! _GENERATED_934 _GENERATED_932 _GENERATED_935 _GENERATED_933 270 285 Filler $T=1790 13860 0 0 $X=1794 $Y=13860
XX30BB92C5137 GND! VDD! _GENERATED_938 _GENERATED_936 _GENERATED_939 _GENERATED_937 271 285 Filler $T=1790 14910 1 0 $X=1794 $Y=14320
XX30BB92C5138 GND! VDD! _GENERATED_942 _GENERATED_940 _GENERATED_943 _GENERATED_941 265 282 Filler $T=2126 9240 0 0 $X=2130 $Y=9240
XX30BB92C5139 GND! VDD! _GENERATED_946 _GENERATED_944 _GENERATED_947 _GENERATED_945 266 282 Filler $T=2126 10290 1 0 $X=2130 $Y=9700
XX30BB92C5140 GND! VDD! _GENERATED_950 _GENERATED_948 _GENERATED_951 _GENERATED_949 266 284 Filler $T=2126 10164 0 0 $X=2130 $Y=10164
XX30BB92C5141 GND! VDD! _GENERATED_954 _GENERATED_952 _GENERATED_955 _GENERATED_953 267 284 Filler $T=2126 11214 1 0 $X=2130 $Y=10624
XX30BB92C5142 GND! VDD! _GENERATED_958 _GENERATED_956 _GENERATED_959 _GENERATED_957 265 280 Filler $T=2126 9366 1 0 $X=2130 $Y=8776
XX30BB92C5143 GND! VDD! _GENERATED_962 _GENERATED_960 _GENERATED_963 _GENERATED_961 272 281 Filler $T=2126 8442 1 0 $X=2130 $Y=7852
XX30BB92C5144 GND! VDD! _GENERATED_966 _GENERATED_964 _GENERATED_967 _GENERATED_965 262 281 Filler $T=2126 7392 0 0 $X=2130 $Y=7392
XX30BB92C5145 GND! VDD! _GENERATED_970 _GENERATED_968 _GENERATED_971 _GENERATED_969 272 280 Filler $T=2126 8316 0 0 $X=2130 $Y=8316
XX30BB92C5146 GND! VDD! _GENERATED_974 _GENERATED_972 _GENERATED_975 _GENERATED_973 268 283 Filler $T=2126 12138 1 0 $X=2130 $Y=11548
XX30BB92C5147 GND! VDD! _GENERATED_978 _GENERATED_976 _GENERATED_979 _GENERATED_977 267 283 Filler $T=2126 11088 0 0 $X=2130 $Y=11088
XX30BB92C5148 GND! VDD! _GENERATED_982 _GENERATED_980 _GENERATED_983 _GENERATED_981 269 287 Filler $T=2126 13062 1 0 $X=2130 $Y=12472
XX30BB92C5149 GND! VDD! _GENERATED_986 _GENERATED_984 _GENERATED_987 _GENERATED_985 268 287 Filler $T=2126 12012 0 0 $X=2130 $Y=12012
XX30BB92C5150 GND! VDD! _GENERATED_990 _GENERATED_988 _GENERATED_991 _GENERATED_989 269 286 Filler $T=2126 12936 0 0 $X=2130 $Y=12936
XX30BB92C5151 GND! VDD! _GENERATED_994 _GENERATED_992 _GENERATED_995 _GENERATED_993 270 286 Filler $T=2126 13986 1 0 $X=2130 $Y=13396
XX30BB92C5152 GND! VDD! _GENERATED_998 _GENERATED_996 _GENERATED_999 _GENERATED_997 270 285 Filler $T=2126 13860 0 0 $X=2130 $Y=13860
XX30BB92C5153 GND! VDD! _GENERATED_1002 _GENERATED_1000 _GENERATED_1003 _GENERATED_1001 271 285 Filler $T=2126 14910 1 0 $X=2130 $Y=14320
XX30BB92C5154 GND! VDD! _GENERATED_1006 _GENERATED_1004 _GENERATED_1007 _GENERATED_1005 271 285 Filler $T=2462 14910 1 0 $X=2466 $Y=14320
XX30BB92C5155 GND! VDD! _GENERATED_1010 _GENERATED_1008 _GENERATED_1011 _GENERATED_1009 270 285 Filler $T=2462 13860 0 0 $X=2466 $Y=13860
XX30BB92C5156 GND! VDD! _GENERATED_1014 _GENERATED_1012 _GENERATED_1015 _GENERATED_1013 270 286 Filler $T=2462 13986 1 0 $X=2466 $Y=13396
XX30BB92C5157 GND! VDD! _GENERATED_1018 _GENERATED_1016 _GENERATED_1019 _GENERATED_1017 269 286 Filler $T=2462 12936 0 0 $X=2466 $Y=12936
XX30BB92C5158 GND! VDD! _GENERATED_1022 _GENERATED_1020 _GENERATED_1023 _GENERATED_1021 268 287 Filler $T=2462 12012 0 0 $X=2466 $Y=12012
XX30BB92C5159 GND! VDD! _GENERATED_1026 _GENERATED_1024 _GENERATED_1027 _GENERATED_1025 269 287 Filler $T=2462 13062 1 0 $X=2466 $Y=12472
XX30BB92C5160 GND! VDD! _GENERATED_1030 _GENERATED_1028 _GENERATED_1031 _GENERATED_1029 267 283 Filler $T=2462 11088 0 0 $X=2466 $Y=11088
XX30BB92C5161 GND! VDD! _GENERATED_1034 _GENERATED_1032 _GENERATED_1035 _GENERATED_1033 268 283 Filler $T=2462 12138 1 0 $X=2466 $Y=11548
XX30BB92C5162 GND! VDD! _GENERATED_1038 _GENERATED_1036 _GENERATED_1039 _GENERATED_1037 267 284 Filler $T=2462 11214 1 0 $X=2466 $Y=10624
XX30BB92C5163 GND! VDD! _GENERATED_1042 _GENERATED_1040 _GENERATED_1043 _GENERATED_1041 266 284 Filler $T=2462 10164 0 0 $X=2466 $Y=10164
XX30BB92C5164 GND! VDD! _GENERATED_1046 _GENERATED_1044 _GENERATED_1047 _GENERATED_1045 266 282 Filler $T=2462 10290 1 0 $X=2466 $Y=9700
XX30BB92C5165 GND! VDD! _GENERATED_1050 _GENERATED_1048 _GENERATED_1051 _GENERATED_1049 265 282 Filler $T=2462 9240 0 0 $X=2466 $Y=9240
XX30BB92C5166 GND! VDD! _GENERATED_1054 _GENERATED_1052 _GENERATED_1055 _GENERATED_1053 265 280 Filler $T=2462 9366 1 0 $X=2466 $Y=8776
XX30BB92C5167 GND! VDD! _GENERATED_1058 _GENERATED_1056 _GENERATED_1059 _GENERATED_1057 272 280 Filler $T=2462 8316 0 0 $X=2466 $Y=8316
XX30BB92C5168 GND! VDD! _GENERATED_1062 _GENERATED_1060 _GENERATED_1063 _GENERATED_1061 272 281 Filler $T=2462 8442 1 0 $X=2466 $Y=7852
XX30BB92C5169 GND! VDD! _GENERATED_1066 _GENERATED_1064 _GENERATED_1067 _GENERATED_1065 262 281 Filler $T=2462 7392 0 0 $X=2466 $Y=7392
XX30BB92C5170 GND! VDD! _GENERATED_1070 _GENERATED_1068 _GENERATED_1071 _GENERATED_1069 271 285 Filler $T=2798 14910 1 0 $X=2802 $Y=14320
XX30BB92C5171 GND! VDD! _GENERATED_1074 _GENERATED_1072 _GENERATED_1075 _GENERATED_1073 270 285 Filler $T=2798 13860 0 0 $X=2802 $Y=13860
XX30BB92C5172 GND! VDD! _GENERATED_1078 _GENERATED_1076 _GENERATED_1079 _GENERATED_1077 270 286 Filler $T=2798 13986 1 0 $X=2802 $Y=13396
XX30BB92C5173 GND! VDD! _GENERATED_1082 _GENERATED_1080 _GENERATED_1083 _GENERATED_1081 269 286 Filler $T=2798 12936 0 0 $X=2802 $Y=12936
XX30BB92C5174 GND! VDD! _GENERATED_1086 _GENERATED_1084 _GENERATED_1087 _GENERATED_1085 268 287 Filler $T=2798 12012 0 0 $X=2802 $Y=12012
XX30BB92C5175 GND! VDD! _GENERATED_1090 _GENERATED_1088 _GENERATED_1091 _GENERATED_1089 269 287 Filler $T=2798 13062 1 0 $X=2802 $Y=12472
XX30BB92C5176 GND! VDD! _GENERATED_1094 _GENERATED_1092 _GENERATED_1095 _GENERATED_1093 267 283 Filler $T=2798 11088 0 0 $X=2802 $Y=11088
XX30BB92C5177 GND! VDD! _GENERATED_1098 _GENERATED_1096 _GENERATED_1099 _GENERATED_1097 268 283 Filler $T=2798 12138 1 0 $X=2802 $Y=11548
XX30BB92C5178 GND! VDD! _GENERATED_1102 _GENERATED_1100 _GENERATED_1103 _GENERATED_1101 272 280 Filler $T=2798 8316 0 0 $X=2802 $Y=8316
XX30BB92C5179 GND! VDD! _GENERATED_1106 _GENERATED_1104 _GENERATED_1107 _GENERATED_1105 262 281 Filler $T=2798 7392 0 0 $X=2802 $Y=7392
XX30BB92C5180 GND! VDD! _GENERATED_1110 _GENERATED_1108 _GENERATED_1111 _GENERATED_1109 272 281 Filler $T=2798 8442 1 0 $X=2802 $Y=7852
XX30BB92C5181 GND! VDD! _GENERATED_1114 _GENERATED_1112 _GENERATED_1115 _GENERATED_1113 265 280 Filler $T=2798 9366 1 0 $X=2802 $Y=8776
XX30BB92C5182 GND! VDD! _GENERATED_1118 _GENERATED_1116 _GENERATED_1119 _GENERATED_1117 267 284 Filler $T=2798 11214 1 0 $X=2802 $Y=10624
XX30BB92C5183 GND! VDD! _GENERATED_1122 _GENERATED_1120 _GENERATED_1123 _GENERATED_1121 266 284 Filler $T=2798 10164 0 0 $X=2802 $Y=10164
XX30BB92C5184 GND! VDD! _GENERATED_1126 _GENERATED_1124 _GENERATED_1127 _GENERATED_1125 266 282 Filler $T=2798 10290 1 0 $X=2802 $Y=9700
XX30BB92C5185 GND! VDD! _GENERATED_1130 _GENERATED_1128 _GENERATED_1131 _GENERATED_1129 265 282 Filler $T=2798 9240 0 0 $X=2802 $Y=9240
XX30BB92C5186 GND! VDD! _GENERATED_1132 VDD! GND! 28 258 278 Filler $T=18874 2898 0 180 $X=18426 $Y=2308
XX30BB92C5187 GND! VDD! GND! _GENERATED_1133 _GENERATED_1134 VDD! 258 275 Filler $T=18422 2772 0 0 $X=18426 $Y=2772
XX30BB92C5188 GND! VDD! GND! _GENERATED_1135 _GENERATED_1136 VDD! 264 VDD! Filler $T=18422 6468 0 0 $X=18426 $Y=6468
XX30BB92C5189 GND! VDD! _GENERATED_1138 VDD! GND! _GENERATED_1137 264 VDD! Filler $T=18874 6594 0 180 $X=18426 $Y=6004
XX30BB92C5190 GND! VDD! GND! _GENERATED_1139 _GENERATED_1140 VDD! 263 VDD! Filler $T=18422 5544 0 0 $X=18426 $Y=5544
XX30BB92C5191 GND! VDD! _GENERATED_1142 VDD! GND! _GENERATED_1141 263 279 Filler $T=18874 5670 0 180 $X=18426 $Y=5080
XX30BB92C5192 GND! VDD! GND! _GENERATED_1143 _GENERATED_1144 VDD! 260 274 Filler $T=18422 3696 0 0 $X=18426 $Y=3696
XX30BB92C5193 GND! VDD! _GENERATED_1146 VDD! GND! _GENERATED_1145 260 275 Filler $T=18874 3822 0 180 $X=18426 $Y=3232
XX30BB92C5194 GND! VDD! _GENERATED_1148 VDD! GND! _GENERATED_1147 261 274 Filler $T=18874 4746 0 180 $X=18426 $Y=4156
XX30BB92C5195 GND! VDD! GND! _GENERATED_1149 _GENERATED_1150 VDD! 261 279 Filler $T=18422 4620 0 0 $X=18426 $Y=4620
XX30BB92C5196 GND! VDD! _GENERATED_1152 VDD! _GENERATED_1153 _GENERATED_1151 262 VDD! Filler $T=9802 7518 0 180 $X=9354 $Y=6928
XX30BB92C5197 GND! VDD! _GENERATED_1156 _GENERATED_1154 _GENERATED_1157 _GENERATED_1155 262 VDD! Filler $T=12826 7518 0 180 $X=12378 $Y=6928
XX30BB92C5198 GND! VDD! _GENERATED_1160 _GENERATED_1158 _GENERATED_1161 _GENERATED_1159 262 VDD! Filler $T=15850 7518 0 180 $X=15402 $Y=6928
XX30BB92C5199 GND! VDD! _GENERATED_1163 VDD! GND! _GENERATED_1162 262 VDD! Filler $T=18874 7518 0 180 $X=18426 $Y=6928
XX30BB92C5200 GND! VDD! Q<3> 94 _GENERATED_1164 273 257 276 tspc_pos_ff $T=17136 0 1 180 $X=15738 $Y=0
XX30BB92C5201 GND! VDD! Q<2> 93 GND! 273 257 276 tspc_pos_ff $T=14112 0 1 180 $X=12714 $Y=0
XX30BB92C5202 GND! VDD! Q<1> 92 GND! 273 257 276 tspc_pos_ff $T=11088 0 1 180 $X=9690 $Y=0
XX30BB92C5203 GND! VDD! Q<0> 91 GND! 273 257 276 tspc_pos_ff $T=8064 0 1 180 $X=6666 $Y=0
XX30BB92C5204 VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! 298 24 
+	23 25 26 27 66 72 73 73 299 300 85 
+	76 90 82 165 166 167 168 86 68 301 100 
+	WS0 302 303 304 261 260 263 264 279 274 275 
+	VDD! VDD! 2to4_decoder_static $T=15738 3234 0 0 $X=15738 $Y=3232
XX30BB92C5205 VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! 305 19 
+	21 20 18 22 65 74 75 75 306 307 85 
+	76 90 82 156 155 154 153 86 68 308 100 
+	WS0 309 310 311 261 260 263 264 279 274 275 
+	VDD! VDD! 2to4_decoder_static $T=12714 3234 0 0 $X=12714 $Y=3232
XX30BB92C5206 VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! 312 9 
+	12 11 10 8 63 77 78 78 313 314 85 
+	76 90 82 132 131 130 129 86 68 315 100 
+	WS0 316 317 318 261 260 263 264 279 274 275 
+	VDD! VDD! 2to4_decoder_static $T=6666 3234 0 0 $X=6666 $Y=3232
XX30BB92C5207 VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 14 
+	13 15 16 17 64 79 80 80 319 320 85 
+	76 90 82 144 143 142 141 86 68 321 100 
+	WS0 322 323 324 261 260 263 264 279 274 275 
+	VDD! VDD! 2to4_decoder_static $T=9690 3234 0 0 $X=9690 $Y=3232
XX30BB92C5208 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=8508 7392 0 0 $X=8508 $Y=7392
XX30BB92C5209 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=7836 7392 0 0 $X=7836 $Y=7392
XX30BB92C5210 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=7164 7392 0 0 $X=7164 $Y=7392
XX30BB92C5211 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=7164 8316 0 0 $X=7164 $Y=8316
XX30BB92C5212 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=7836 8316 0 0 $X=7836 $Y=8316
XX30BB92C5213 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=8508 8316 0 0 $X=8508 $Y=8316
XX30BB92C5214 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=9180 8316 0 0 $X=9180 $Y=8316
XX30BB92C5215 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=9180 7392 0 0 $X=9180 $Y=7392
XX30BB92C5216 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=9180 9240 0 0 $X=9180 $Y=9240
XX30BB92C5217 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=7164 9240 0 0 $X=7164 $Y=9240
XX30BB92C5218 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=7836 9240 0 0 $X=7836 $Y=9240
XX30BB92C5219 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=8508 9240 0 0 $X=8508 $Y=9240
XX30BB92C5220 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=9180 10164 0 0 $X=9180 $Y=10164
XX30BB92C5221 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=8508 10164 0 0 $X=8508 $Y=10164
XX30BB92C5222 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=7836 10164 0 0 $X=7836 $Y=10164
XX30BB92C5223 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=7164 10164 0 0 $X=7164 $Y=10164
XX30BB92C5224 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=8508 11088 0 0 $X=8508 $Y=11088
XX30BB92C5225 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=7836 11088 0 0 $X=7836 $Y=11088
XX30BB92C5226 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=7164 11088 0 0 $X=7164 $Y=11088
XX30BB92C5227 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=9180 11088 0 0 $X=9180 $Y=11088
XX30BB92C5228 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=7164 12012 0 0 $X=7164 $Y=12012
XX30BB92C5229 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=7836 12012 0 0 $X=7836 $Y=12012
XX30BB92C5230 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=8508 12012 0 0 $X=8508 $Y=12012
XX30BB92C5231 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=9180 12012 0 0 $X=9180 $Y=12012
XX30BB92C5232 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=9180 12936 0 0 $X=9180 $Y=12936
XX30BB92C5233 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=7164 12936 0 0 $X=7164 $Y=12936
XX30BB92C5234 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=7836 12936 0 0 $X=7836 $Y=12936
XX30BB92C5235 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=8508 12936 0 0 $X=8508 $Y=12936
XX30BB92C5236 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=9180 13860 0 0 $X=9180 $Y=13860
XX30BB92C5237 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=8508 13860 0 0 $X=8508 $Y=13860
XX30BB92C5238 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=7836 13860 0 0 $X=7836 $Y=13860
XX30BB92C5239 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=7164 13860 0 0 $X=7164 $Y=13860
XX30BB92C5240 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=10188 13860 0 0 $X=10188 $Y=13860
XX30BB92C5241 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=10860 13860 0 0 $X=10860 $Y=13860
XX30BB92C5242 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=11532 13860 0 0 $X=11532 $Y=13860
XX30BB92C5243 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=12204 13860 0 0 $X=12204 $Y=13860
XX30BB92C5244 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=11532 12936 0 0 $X=11532 $Y=12936
XX30BB92C5245 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=10860 12936 0 0 $X=10860 $Y=12936
XX30BB92C5246 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=10188 12936 0 0 $X=10188 $Y=12936
XX30BB92C5247 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=12204 12936 0 0 $X=12204 $Y=12936
XX30BB92C5248 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=12204 12012 0 0 $X=12204 $Y=12012
XX30BB92C5249 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=11532 12012 0 0 $X=11532 $Y=12012
XX30BB92C5250 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=10860 12012 0 0 $X=10860 $Y=12012
XX30BB92C5251 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=10188 12012 0 0 $X=10188 $Y=12012
XX30BB92C5252 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=12204 11088 0 0 $X=12204 $Y=11088
XX30BB92C5253 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=10188 11088 0 0 $X=10188 $Y=11088
XX30BB92C5254 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=10860 11088 0 0 $X=10860 $Y=11088
XX30BB92C5255 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=11532 11088 0 0 $X=11532 $Y=11088
XX30BB92C5256 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=10188 10164 0 0 $X=10188 $Y=10164
XX30BB92C5257 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=10860 10164 0 0 $X=10860 $Y=10164
XX30BB92C5258 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=11532 10164 0 0 $X=11532 $Y=10164
XX30BB92C5259 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=12204 10164 0 0 $X=12204 $Y=10164
XX30BB92C5260 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=11532 9240 0 0 $X=11532 $Y=9240
XX30BB92C5261 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=10860 9240 0 0 $X=10860 $Y=9240
XX30BB92C5262 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=10188 9240 0 0 $X=10188 $Y=9240
XX30BB92C5263 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=12204 9240 0 0 $X=12204 $Y=9240
XX30BB92C5264 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=10188 8316 0 0 $X=10188 $Y=8316
XX30BB92C5265 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=10860 8316 0 0 $X=10860 $Y=8316
XX30BB92C5266 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=11532 8316 0 0 $X=11532 $Y=8316
XX30BB92C5267 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=12204 8316 0 0 $X=12204 $Y=8316
XX30BB92C5268 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=12204 7392 0 0 $X=12204 $Y=7392
XX30BB92C5269 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=11532 7392 0 0 $X=11532 $Y=7392
XX30BB92C5270 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=10188 7392 0 0 $X=10188 $Y=7392
XX30BB92C5271 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=10860 7392 0 0 $X=10860 $Y=7392
XX30BB92C5272 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=18252 9240 0 0 $X=18252 $Y=9240
XX30BB92C5273 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=16236 9240 0 0 $X=16236 $Y=9240
XX30BB92C5274 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=16908 9240 0 0 $X=16908 $Y=9240
XX30BB92C5275 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=17580 9240 0 0 $X=17580 $Y=9240
XX30BB92C5276 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=18252 10164 0 0 $X=18252 $Y=10164
XX30BB92C5277 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=17580 10164 0 0 $X=17580 $Y=10164
XX30BB92C5278 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=16908 10164 0 0 $X=16908 $Y=10164
XX30BB92C5279 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=16236 10164 0 0 $X=16236 $Y=10164
XX30BB92C5280 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=17580 11088 0 0 $X=17580 $Y=11088
XX30BB92C5281 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=16908 11088 0 0 $X=16908 $Y=11088
XX30BB92C5282 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=16236 11088 0 0 $X=16236 $Y=11088
XX30BB92C5283 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=18252 11088 0 0 $X=18252 $Y=11088
XX30BB92C5284 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=16236 12012 0 0 $X=16236 $Y=12012
XX30BB92C5285 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=16908 12012 0 0 $X=16908 $Y=12012
XX30BB92C5286 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=17580 12012 0 0 $X=17580 $Y=12012
XX30BB92C5287 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=18252 12012 0 0 $X=18252 $Y=12012
XX30BB92C5288 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=18252 12936 0 0 $X=18252 $Y=12936
XX30BB92C5289 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=16236 12936 0 0 $X=16236 $Y=12936
XX30BB92C5290 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=16908 12936 0 0 $X=16908 $Y=12936
XX30BB92C5291 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=17580 12936 0 0 $X=17580 $Y=12936
XX30BB92C5292 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=18252 13860 0 0 $X=18252 $Y=13860
XX30BB92C5293 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=17580 13860 0 0 $X=17580 $Y=13860
XX30BB92C5294 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=16908 13860 0 0 $X=16908 $Y=13860
XX30BB92C5295 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=16236 13860 0 0 $X=16236 $Y=13860
XX30BB92C5296 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=14556 13860 0 0 $X=14556 $Y=13860
XX30BB92C5297 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=15228 13860 0 0 $X=15228 $Y=13860
XX30BB92C5298 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=14556 12936 0 0 $X=14556 $Y=12936
XX30BB92C5299 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=15228 12936 0 0 $X=15228 $Y=12936
XX30BB92C5300 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=15228 12012 0 0 $X=15228 $Y=12012
XX30BB92C5301 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=14556 12012 0 0 $X=14556 $Y=12012
XX30BB92C5302 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=15228 11088 0 0 $X=15228 $Y=11088
XX30BB92C5303 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=14556 11088 0 0 $X=14556 $Y=11088
XX30BB92C5304 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=14556 10164 0 0 $X=14556 $Y=10164
XX30BB92C5305 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=15228 10164 0 0 $X=15228 $Y=10164
XX30BB92C5306 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=14556 9240 0 0 $X=14556 $Y=9240
XX30BB92C5307 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=15228 9240 0 0 $X=15228 $Y=9240
XX30BB92C5308 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=16908 7392 0 0 $X=16908 $Y=7392
XX30BB92C5309 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=16236 7392 0 0 $X=16236 $Y=7392
XX30BB92C5310 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=17580 7392 0 0 $X=17580 $Y=7392
XX30BB92C5311 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=18252 7392 0 0 $X=18252 $Y=7392
XX30BB92C5312 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=18252 8316 0 0 $X=18252 $Y=8316
XX30BB92C5313 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=17580 8316 0 0 $X=17580 $Y=8316
XX30BB92C5314 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=16908 8316 0 0 $X=16908 $Y=8316
XX30BB92C5315 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=16236 8316 0 0 $X=16236 $Y=8316
XX30BB92C5316 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=13212 13860 0 0 $X=13212 $Y=13860
XX30BB92C5317 GND! VDD! GND! 270 271 285 bitcell_precharge_filler $T=13884 13860 0 0 $X=13884 $Y=13860
XX30BB92C5318 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=13884 12936 0 0 $X=13884 $Y=12936
XX30BB92C5319 GND! VDD! GND! 269 270 286 bitcell_precharge_filler $T=13212 12936 0 0 $X=13212 $Y=12936
XX30BB92C5320 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=13884 12012 0 0 $X=13884 $Y=12012
XX30BB92C5321 GND! VDD! GND! 268 269 287 bitcell_precharge_filler $T=13212 12012 0 0 $X=13212 $Y=12012
XX30BB92C5322 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=13212 11088 0 0 $X=13212 $Y=11088
XX30BB92C5323 GND! VDD! GND! 267 268 283 bitcell_precharge_filler $T=13884 11088 0 0 $X=13884 $Y=11088
XX30BB92C5324 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=13212 10164 0 0 $X=13212 $Y=10164
XX30BB92C5325 GND! VDD! GND! 266 267 284 bitcell_precharge_filler $T=13884 10164 0 0 $X=13884 $Y=10164
XX30BB92C5326 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=13884 9240 0 0 $X=13884 $Y=9240
XX30BB92C5327 GND! VDD! GND! 265 266 282 bitcell_precharge_filler $T=13212 9240 0 0 $X=13212 $Y=9240
XX30BB92C5328 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=13212 8316 0 0 $X=13212 $Y=8316
XX30BB92C5329 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=13884 8316 0 0 $X=13884 $Y=8316
XX30BB92C5330 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=14556 8316 0 0 $X=14556 $Y=8316
XX30BB92C5331 GND! VDD! GND! 272 265 280 bitcell_precharge_filler $T=15228 8316 0 0 $X=15228 $Y=8316
XX30BB92C5332 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=15228 7392 0 0 $X=15228 $Y=7392
XX30BB92C5333 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=14556 7392 0 0 $X=14556 $Y=7392
XX30BB92C5334 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=13212 7392 0 0 $X=13212 $Y=7392
XX30BB92C5335 GND! VDD! GND! 262 272 281 bitcell_precharge_filler $T=13884 7392 0 0 $X=13884 $Y=7392
XX30BB92C5336 VDD! GND! GND! GND! VDD! VDD! GND! VDD! GND! GND! VDD! 
+	GND! VDD! GND! GND! VDD! 511 A<2> A<3> 508 A<4> 485 
+	96 104 99 105 106 98 103 108 107 262 272 
+	266 265 268 267 271 270 269 281 280 282 284 
+	283 286 287 285 486 484 static_row_decoder_3by8 $T=2486 13270 0 0 $X=3138 $Y=7391
XX30BB92C5337 GND! VDD! VDD! GND! 257 276 2to4_decoder_static_filler_17 $T=18870 1054 0 180 $X=18426 $Y=462
XX30BB92C5338 GND! VDD! _GENERATED_1166 _GENERATED_1165 257 277 2to4_decoder_static_filler_17 $T=18426 920 0 0 $X=18426 $Y=924
XX30BB92C5339 GND! VDD! _GENERATED_1168 _GENERATED_1167 257 277 2to4_decoder_static_filler_17 $T=17754 920 0 0 $X=17754 $Y=924
XX30BB92C5340 GND! VDD! _GENERATED_1170 _GENERATED_1169 257 277 2to4_decoder_static_filler_17 $T=18090 920 0 0 $X=18090 $Y=924
XX30BB92C5341 GND! VDD! _GENERATED_1172 _GENERATED_1171 257 276 2to4_decoder_static_filler_17 $T=18534 1054 0 180 $X=18090 $Y=462
XX30BB92C5342 GND! VDD! _GENERATED_1174 _GENERATED_1173 257 276 2to4_decoder_static_filler_17 $T=18198 1054 0 180 $X=17754 $Y=462
XX30BB92C5343 GND! VDD! _GENERATED_1176 _GENERATED_1175 257 276 2to4_decoder_static_filler_17 $T=17526 1054 0 180 $X=17082 $Y=462
XX30BB92C5344 GND! VDD! _GENERATED_1178 _GENERATED_1177 257 276 2to4_decoder_static_filler_17 $T=17862 1054 0 180 $X=17418 $Y=462
XX30BB92C5345 GND! VDD! _GENERATED_1180 _GENERATED_1179 257 277 2to4_decoder_static_filler_17 $T=14730 920 0 0 $X=14730 $Y=924
XX30BB92C5346 GND! VDD! _GENERATED_1182 _GENERATED_1181 257 277 2to4_decoder_static_filler_17 $T=15066 920 0 0 $X=15066 $Y=924
XX30BB92C5347 GND! VDD! _GENERATED_1184 _GENERATED_1183 257 277 2to4_decoder_static_filler_17 $T=15402 920 0 0 $X=15402 $Y=924
XX30BB92C5348 GND! VDD! _GENERATED_1186 _GENERATED_1185 257 276 2to4_decoder_static_filler_17 $T=15846 1054 0 180 $X=15402 $Y=462
XX30BB92C5349 GND! VDD! _GENERATED_1188 _GENERATED_1187 257 276 2to4_decoder_static_filler_17 $T=15510 1054 0 180 $X=15065 $Y=462
XX30BB92C5350 GND! VDD! _GENERATED_1190 _GENERATED_1189 257 276 2to4_decoder_static_filler_17 $T=15174 1054 0 180 $X=14729 $Y=462
XX30BB92C5351 GND! VDD! _GENERATED_1192 _GENERATED_1191 257 276 2to4_decoder_static_filler_17 $T=14838 1054 0 180 $X=14394 $Y=462
XX30BB92C5352 GND! VDD! _GENERATED_1194 _GENERATED_1193 257 276 2to4_decoder_static_filler_17 $T=14502 1054 0 180 $X=14058 $Y=462
XX30BB92C5353 GND! VDD! _GENERATED_1196 _GENERATED_1195 257 276 2to4_decoder_static_filler_17 $T=11814 1054 0 180 $X=11370 $Y=462
XX30BB92C5354 GND! VDD! _GENERATED_1198 _GENERATED_1197 257 276 2to4_decoder_static_filler_17 $T=11478 1054 0 180 $X=11033 $Y=462
XX30BB92C5355 GND! VDD! _GENERATED_1200 _GENERATED_1199 257 276 2to4_decoder_static_filler_17 $T=12150 1054 0 180 $X=11706 $Y=462
XX30BB92C5356 GND! VDD! _GENERATED_1202 _GENERATED_1201 257 276 2to4_decoder_static_filler_17 $T=12486 1054 0 180 $X=12042 $Y=462
XX30BB92C5357 GND! VDD! _GENERATED_1204 _GENERATED_1203 257 277 2to4_decoder_static_filler_17 $T=12042 920 0 0 $X=12042 $Y=924
XX30BB92C5358 GND! VDD! _GENERATED_1206 _GENERATED_1205 257 277 2to4_decoder_static_filler_17 $T=11706 920 0 0 $X=11706 $Y=924
XX30BB92C5359 GND! VDD! _GENERATED_1208 _GENERATED_1207 257 277 2to4_decoder_static_filler_17 $T=12378 920 0 0 $X=12378 $Y=924
XX30BB92C5360 GND! VDD! _GENERATED_1210 _GENERATED_1209 257 276 2to4_decoder_static_filler_17 $T=12822 1054 0 180 $X=12378 $Y=462
XX30BB92C5361 GND! VDD! _GENERATED_1212 _GENERATED_1211 257 276 2to4_decoder_static_filler_17 $T=8454 1054 0 180 $X=8010 $Y=462
XX30BB92C5362 GND! VDD! _GENERATED_1214 _GENERATED_1213 257 276 2to4_decoder_static_filler_17 $T=8790 1054 0 180 $X=8346 $Y=462
XX30BB92C5363 GND! VDD! _GENERATED_1216 _GENERATED_1215 257 276 2to4_decoder_static_filler_17 $T=9126 1054 0 180 $X=8681 $Y=462
XX30BB92C5364 GND! VDD! _GENERATED_1218 _GENERATED_1217 257 276 2to4_decoder_static_filler_17 $T=9462 1054 0 180 $X=9017 $Y=462
XX30BB92C5365 GND! VDD! _GENERATED_1220 _GENERATED_1219 257 276 2to4_decoder_static_filler_17 $T=9798 1054 0 180 $X=9354 $Y=462
XX30BB92C5366 GND! VDD! _GENERATED_1222 _GENERATED_1221 257 277 2to4_decoder_static_filler_17 $T=9354 920 0 0 $X=9354 $Y=924
XX30BB92C5367 GND! VDD! _GENERATED_1224 _GENERATED_1223 257 277 2to4_decoder_static_filler_17 $T=9018 920 0 0 $X=9018 $Y=924
XX30BB92C5368 GND! VDD! _GENERATED_1226 _GENERATED_1225 257 277 2to4_decoder_static_filler_17 $T=8682 920 0 0 $X=8682 $Y=924
XX30BB92C5369 GND! VDD! 73 338 24 127 94 D<3> D<3> 126 128 
+	128 257 277 483 read_circuit $T=15738 920 0 0 $X=15738 $Y=924
XX30BB92C5370 GND! VDD! 75 339 19 124 93 D<2> D<2> 123 125 
+	125 257 277 481 read_circuit $T=12714 920 0 0 $X=12714 $Y=924
XX30BB92C5371 GND! VDD! 80 340 14 121 92 D<1> D<1> 120 122 
+	122 257 277 482 read_circuit $T=9690 920 0 0 $X=9690 $Y=924
XX30BB92C5372 GND! VDD! 78 328 9 118 91 D<0> D<0> 117 119 
+	119 257 277 480 read_circuit $T=6666 920 0 0 $X=6666 $Y=924
XX30BB92C5373 GND! VDD! _GENERATED_1228 _GENERATED_1227 273 276 sram_filler $T=18422 0 0 0 $X=18426 $Y=0
XX30BB92C5374 GND! VDD! _GENERATED_1230 _GENERATED_1229 273 276 sram_filler $T=17078 0 0 0 $X=17082 $Y=0
XX30BB92C5375 GND! VDD! _GENERATED_1232 _GENERATED_1231 273 276 sram_filler $T=17414 0 0 0 $X=17418 $Y=0
XX30BB92C5376 GND! VDD! _GENERATED_1234 _GENERATED_1233 273 276 sram_filler $T=17750 0 0 0 $X=17754 $Y=0
XX30BB92C5377 GND! VDD! _GENERATED_1236 _GENERATED_1235 273 276 sram_filler $T=18086 0 0 0 $X=18090 $Y=0
XX30BB92C5378 GND! VDD! _GENERATED_1238 _GENERATED_1237 273 276 sram_filler $T=15398 0 0 0 $X=15402 $Y=0
XX30BB92C5379 GND! VDD! _GENERATED_1240 _GENERATED_1239 273 276 sram_filler $T=15062 0 0 0 $X=15066 $Y=0
XX30BB92C5380 GND! VDD! _GENERATED_1242 _GENERATED_1241 273 276 sram_filler $T=14726 0 0 0 $X=14730 $Y=0
XX30BB92C5381 GND! VDD! _GENERATED_1244 _GENERATED_1243 273 276 sram_filler $T=6326 0 0 0 $X=6330 $Y=0
XX30BB92C5382 GND! VDD! _GENERATED_1246 _GENERATED_1245 273 276 sram_filler $T=5990 0 0 0 $X=5994 $Y=0
XX30BB92C5383 GND! VDD! _GENERATED_1248 _GENERATED_1247 273 276 sram_filler $T=5654 0 0 0 $X=5657 $Y=0
XX30BB92C5384 GND! VDD! _GENERATED_1250 _GENERATED_1249 273 276 sram_filler $T=5318 0 0 0 $X=5322 $Y=0
XX30BB92C5385 GND! VDD! _GENERATED_1252 _GENERATED_1251 273 276 sram_filler $T=8006 0 0 0 $X=8010 $Y=0
XX30BB92C5386 GND! VDD! _GENERATED_1254 _GENERATED_1253 273 276 sram_filler $T=8342 0 0 0 $X=8346 $Y=0
XX30BB92C5387 GND! VDD! _GENERATED_1256 _GENERATED_1255 273 276 sram_filler $T=8678 0 0 0 $X=8682 $Y=0
XX30BB92C5388 GND! VDD! _GENERATED_1258 _GENERATED_1257 273 276 sram_filler $T=14054 0 0 0 $X=14058 $Y=0
XX30BB92C5389 GND! VDD! _GENERATED_1260 _GENERATED_1259 273 276 sram_filler $T=12038 0 0 0 $X=12042 $Y=0
XX30BB92C5390 GND! VDD! _GENERATED_1262 _GENERATED_1261 273 276 sram_filler $T=11702 0 0 0 $X=11706 $Y=0
XX30BB92C5391 GND! VDD! _GENERATED_1264 _GENERATED_1263 273 276 sram_filler $T=11366 0 0 0 $X=11370 $Y=0
XX30BB92C5392 GND! VDD! _GENERATED_1266 _GENERATED_1265 273 276 sram_filler $T=11030 0 0 0 $X=11033 $Y=0
XX30BB92C5393 GND! VDD! _GENERATED_1268 _GENERATED_1267 273 276 sram_filler $T=14390 0 0 0 $X=14394 $Y=0
XX30BB92C5394 GND! VDD! _GENERATED_1270 _GENERATED_1269 273 276 sram_filler $T=9014 0 0 0 $X=9017 $Y=0
XX30BB92C5395 GND! VDD! _GENERATED_1272 _GENERATED_1271 273 276 sram_filler $T=9350 0 0 0 $X=9354 $Y=0
XX30BB92C5396 GND! VDD! _GENERATED_1274 _GENERATED_1273 273 276 sram_filler $T=12374 0 0 0 $X=12378 $Y=0
XX30BB92C5397 GND! VDD! _GENERATED_1276 _GENERATED_1275 273 276 sram_filler $T=4982 0 0 0 $X=4986 $Y=0
XX30BB92C5398 GND! VDD! _GENERATED_1278 _GENERATED_1277 273 276 sram_filler $T=4646 0 0 0 $X=4649 $Y=0
XX30BB92C5399 GND! VDD! _GENERATED_1280 _GENERATED_1279 273 276 sram_filler $T=4310 0 0 0 $X=4314 $Y=0
XX30BB92C5400 GND! VDD! _GENERATED_1282 _GENERATED_1281 273 276 sram_filler $T=3974 0 0 0 $X=3978 $Y=0
XX30BB92C5401 GND! VDD! _GENERATED_1284 _GENERATED_1283 273 276 sram_filler $T=2630 0 0 0 $X=2634 $Y=0
XX30BB92C5402 GND! VDD! _GENERATED_1286 _GENERATED_1285 273 276 sram_filler $T=2966 0 0 0 $X=2970 $Y=0
XX30BB92C5403 GND! VDD! _GENERATED_1288 _GENERATED_1287 273 276 sram_filler $T=3302 0 0 0 $X=3306 $Y=0
XX30BB92C5404 GND! VDD! _GENERATED_1290 _GENERATED_1289 273 276 sram_filler $T=3638 0 0 0 $X=3642 $Y=0
XX30BB92C5405 GND! VDD! _GENERATED_1292 _GENERATED_1291 273 276 sram_filler $T=1286 0 0 0 $X=1290 $Y=0
XX30BB92C5406 GND! VDD! _GENERATED_1294 _GENERATED_1293 273 276 sram_filler $T=1622 0 0 0 $X=1626 $Y=0
XX30BB92C5407 GND! VDD! _GENERATED_1296 _GENERATED_1295 273 276 sram_filler $T=1958 0 0 0 $X=1962 $Y=0
XX30BB92C5408 GND! VDD! _GENERATED_1298 _GENERATED_1297 273 276 sram_filler $T=2294 0 0 0 $X=2298 $Y=0
XX30BB92C5409 GND! VDD! _GENERATED_1300 _GENERATED_1299 273 276 sram_filler $T=950 0 0 0 $X=954 $Y=0
XX30BB92C5410 GND! VDD! _GENERATED_1302 _GENERATED_1301 273 276 sram_filler $T=614 0 0 0 $X=618 $Y=0
XX30BB92C5411 GND! VDD! _GENERATED_1304 _GENERATED_1303 273 276 sram_filler $T=278 0 0 0 $X=282 $Y=0
XX30BB92C5412 GND! VDD! _GENERATED_1306 _GENERATED_1305 273 276 sram_filler $T=-58 0 0 0 $X=-54 $Y=0
XX30BB92C5413 GND! VDD! _GENERATED_1308 _GENERATED_1307 257 277 sram_filler $T=950 924 0 0 $X=954 $Y=924
XX30BB92C5414 GND! VDD! _GENERATED_1310 _GENERATED_1309 257 277 sram_filler $T=614 924 0 0 $X=618 $Y=924
XX30BB92C5415 GND! VDD! _GENERATED_1312 _GENERATED_1311 257 277 sram_filler $T=278 924 0 0 $X=282 $Y=924
XX30BB92C5416 GND! VDD! _GENERATED_1314 _GENERATED_1313 257 277 sram_filler $T=-58 924 0 0 $X=-54 $Y=924
XX30BB92C5417 GND! VDD! _GENERATED_1316 _GENERATED_1315 259 278 sram_filler $T=950 1848 0 0 $X=954 $Y=1848
XX30BB92C5418 GND! VDD! _GENERATED_1318 _GENERATED_1317 259 278 sram_filler $T=614 1848 0 0 $X=618 $Y=1848
XX30BB92C5419 GND! VDD! _GENERATED_1320 _GENERATED_1319 259 278 sram_filler $T=278 1848 0 0 $X=282 $Y=1848
XX30BB92C5420 GND! VDD! _GENERATED_1322 _GENERATED_1321 259 278 sram_filler $T=-58 1848 0 0 $X=-54 $Y=1848
XX30BB92C5421 GND! VDD! _GENERATED_1324 _GENERATED_1323 258 275 sram_filler $T=-58 2772 0 0 $X=-54 $Y=2772
XX30BB92C5422 GND! VDD! _GENERATED_1326 _GENERATED_1325 258 275 sram_filler $T=278 2772 0 0 $X=282 $Y=2772
XX30BB92C5423 GND! VDD! _GENERATED_1328 _GENERATED_1327 258 275 sram_filler $T=614 2772 0 0 $X=618 $Y=2772
XX30BB92C5424 GND! VDD! _GENERATED_1330 _GENERATED_1329 258 275 sram_filler $T=950 2772 0 0 $X=954 $Y=2772
XX30BB92C5425 GND! VDD! _GENERATED_1332 _GENERATED_1331 260 274 sram_filler $T=-58 3696 0 0 $X=-54 $Y=3696
XX30BB92C5426 GND! VDD! _GENERATED_1334 _GENERATED_1333 260 274 sram_filler $T=278 3696 0 0 $X=282 $Y=3696
XX30BB92C5427 GND! VDD! _GENERATED_1336 _GENERATED_1335 260 274 sram_filler $T=614 3696 0 0 $X=618 $Y=3696
XX30BB92C5428 GND! VDD! _GENERATED_1338 _GENERATED_1337 260 274 sram_filler $T=950 3696 0 0 $X=954 $Y=3696
XX30BB92C5429 GND! VDD! VDD! _GENERATED_1339 259 278 sram_filler $T=6326 1848 0 0 $X=6330 $Y=1848
XX30BB92C5430 GND! VDD! _GENERATED_1341 _GENERATED_1340 259 278 sram_filler $T=5486 1848 0 0 $X=5489 $Y=1848
XX30BB92C5431 GND! VDD! _GENERATED_1343 _GENERATED_1342 259 278 sram_filler $T=5822 1848 0 0 $X=5826 $Y=1848
XX30BB92C5432 GND! VDD! _GENERATED_1344 GND! 259 278 sram_filler $T=6158 1848 0 0 $X=6162 $Y=1848
XX30BB92C5433 GND! VDD! VDD! _GENERATED_1345 258 275 sram_filler $T=18086 2772 0 0 $X=18090 $Y=2772
XX30BB92C5434 GND! VDD! _GENERATED_1347 _GENERATED_1346 258 275 sram_filler $T=17582 2772 0 0 $X=17586 $Y=2772
XX30BB92C5435 GND! VDD! _GENERATED_1348 GND! 258 275 sram_filler $T=17918 2772 0 0 $X=17922 $Y=2772
XX30BB92C5436 GND! VDD! _GENERATED_1350 _GENERATED_1349 258 275 sram_filler $T=17246 2772 0 0 $X=17250 $Y=2772
XX30BB92C5437 GND! VDD! _GENERATED_1352 _GENERATED_1351 258 275 sram_filler $T=16910 2772 0 0 $X=16914 $Y=2772
XX30BB92C5438 GND! VDD! _GENERATED_1354 _GENERATED_1353 258 275 sram_filler $T=16238 2772 0 0 $X=16242 $Y=2772
XX30BB92C5439 GND! VDD! _GENERATED_1356 _GENERATED_1355 258 275 sram_filler $T=16574 2772 0 0 $X=16578 $Y=2772
XX30BB92C5440 GND! VDD! _GENERATED_1358 _GENERATED_1357 258 275 sram_filler $T=13550 2772 0 0 $X=13554 $Y=2772
XX30BB92C5441 GND! VDD! _GENERATED_1360 _GENERATED_1359 258 275 sram_filler $T=12878 2772 0 0 $X=12882 $Y=2772
XX30BB92C5442 GND! VDD! _GENERATED_1362 _GENERATED_1361 258 275 sram_filler $T=13214 2772 0 0 $X=13218 $Y=2772
XX30BB92C5443 GND! VDD! _GENERATED_1364 _GENERATED_1363 258 275 sram_filler $T=12542 2772 0 0 $X=12546 $Y=2772
XX30BB92C5444 GND! VDD! _GENERATED_1366 _GENERATED_1365 258 275 sram_filler $T=12206 2772 0 0 $X=12209 $Y=2772
XX30BB92C5445 GND! VDD! _GENERATED_1368 _GENERATED_1367 258 275 sram_filler $T=11534 2772 0 0 $X=11538 $Y=2772
XX30BB92C5446 GND! VDD! _GENERATED_1370 _GENERATED_1369 258 275 sram_filler $T=11870 2772 0 0 $X=11874 $Y=2772
XX30BB92C5447 GND! VDD! _GENERATED_1372 _GENERATED_1371 258 275 sram_filler $T=11198 2772 0 0 $X=11202 $Y=2772
XX30BB92C5448 GND! VDD! _GENERATED_1374 _GENERATED_1373 258 275 sram_filler $T=10862 2772 0 0 $X=10866 $Y=2772
XX30BB92C5449 GND! VDD! _GENERATED_1376 _GENERATED_1375 258 275 sram_filler $T=15566 2772 0 0 $X=15570 $Y=2772
XX30BB92C5450 GND! VDD! _GENERATED_1378 _GENERATED_1377 258 275 sram_filler $T=15902 2772 0 0 $X=15906 $Y=2772
XX30BB92C5451 GND! VDD! _GENERATED_1380 _GENERATED_1379 258 275 sram_filler $T=15230 2772 0 0 $X=15234 $Y=2772
XX30BB92C5452 GND! VDD! _GENERATED_1382 _GENERATED_1381 258 275 sram_filler $T=14894 2772 0 0 $X=14898 $Y=2772
XX30BB92C5453 GND! VDD! _GENERATED_1384 _GENERATED_1383 258 275 sram_filler $T=14222 2772 0 0 $X=14226 $Y=2772
XX30BB92C5454 GND! VDD! _GENERATED_1386 _GENERATED_1385 258 275 sram_filler $T=14558 2772 0 0 $X=14562 $Y=2772
XX30BB92C5455 GND! VDD! _GENERATED_1388 _GENERATED_1387 258 275 sram_filler $T=13886 2772 0 0 $X=13890 $Y=2772
XX30BB92C5456 GND! VDD! _GENERATED_1390 _GENERATED_1389 258 275 sram_filler $T=10190 2772 0 0 $X=10193 $Y=2772
XX30BB92C5457 GND! VDD! _GENERATED_1392 _GENERATED_1391 258 275 sram_filler $T=10526 2772 0 0 $X=10530 $Y=2772
XX30BB92C5458 GND! VDD! _GENERATED_1394 _GENERATED_1393 258 275 sram_filler $T=9854 2772 0 0 $X=9858 $Y=2772
XX30BB92C5459 GND! VDD! _GENERATED_1396 _GENERATED_1395 258 275 sram_filler $T=9518 2772 0 0 $X=9522 $Y=2772
XX30BB92C5460 GND! VDD! _GENERATED_1398 _GENERATED_1397 258 275 sram_filler $T=8846 2772 0 0 $X=8850 $Y=2772
XX30BB92C5461 GND! VDD! _GENERATED_1400 _GENERATED_1399 258 275 sram_filler $T=9182 2772 0 0 $X=9186 $Y=2772
XX30BB92C5462 GND! VDD! _GENERATED_1402 _GENERATED_1401 258 275 sram_filler $T=8510 2772 0 0 $X=8514 $Y=2772
XX30BB92C5463 GND! VDD! _GENERATED_1404 _GENERATED_1403 258 275 sram_filler $T=8174 2772 0 0 $X=8177 $Y=2772
XX30BB92C5464 GND! VDD! _GENERATED_1406 _GENERATED_1405 258 275 sram_filler $T=7502 2772 0 0 $X=7505 $Y=2772
XX30BB92C5465 GND! VDD! _GENERATED_1408 _GENERATED_1407 258 275 sram_filler $T=7838 2772 0 0 $X=7842 $Y=2772
XX30BB92C5466 GND! VDD! _GENERATED_1410 _GENERATED_1409 258 275 sram_filler $T=7166 2772 0 0 $X=7170 $Y=2772
XX30BB92C5467 GND! VDD! _GENERATED_1412 _GENERATED_1411 258 275 sram_filler $T=6830 2772 0 0 $X=6834 $Y=2772
XX30BB92C5468 GND! VDD! _GENERATED_1414 _GENERATED_1413 258 275 sram_filler $T=6158 2772 0 0 $X=6162 $Y=2772
XX30BB92C5469 GND! VDD! _GENERATED_1416 _GENERATED_1415 258 275 sram_filler $T=6494 2772 0 0 $X=6497 $Y=2772
XX30BB92C5470 GND! VDD! _GENERATED_1418 _GENERATED_1417 258 275 sram_filler $T=5822 2772 0 0 $X=5826 $Y=2772
XX30BB92C5471 GND! VDD! _GENERATED_1420 _GENERATED_1419 258 275 sram_filler $T=5486 2772 0 0 $X=5489 $Y=2772
XX30BB92C5472 GND! VDD! _GENERATED_1422 _GENERATED_1421 264 VDD! sram_filler $T=15398 6468 0 0 $X=15402 $Y=6468
XX30BB92C5473 GND! VDD! _GENERATED_1424 _GENERATED_1423 263 VDD! sram_filler $T=15398 5544 0 0 $X=15402 $Y=5544
XX30BB92C5474 GND! VDD! _GENERATED_1426 _GENERATED_1425 261 279 sram_filler $T=15398 4620 0 0 $X=15402 $Y=4620
XX30BB92C5475 GND! VDD! _GENERATED_1428 _GENERATED_1427 260 274 sram_filler $T=15398 3696 0 0 $X=15402 $Y=3696
XX30BB92C5476 GND! VDD! _GENERATED_1430 _GENERATED_1429 261 279 sram_filler $T=12374 4620 0 0 $X=12378 $Y=4620
XX30BB92C5477 GND! VDD! _GENERATED_1432 _GENERATED_1431 260 274 sram_filler $T=12374 3696 0 0 $X=12378 $Y=3696
XX30BB92C5478 GND! VDD! _GENERATED_1434 _GENERATED_1433 263 VDD! sram_filler $T=12374 5544 0 0 $X=12378 $Y=5544
XX30BB92C5479 GND! VDD! _GENERATED_1436 _GENERATED_1435 264 VDD! sram_filler $T=12374 6468 0 0 $X=12378 $Y=6468
XX30BB92C5480 GND! VDD! _GENERATED_1438 _GENERATED_1437 260 274 sram_filler $T=9350 3696 0 0 $X=9354 $Y=3696
XX30BB92C5481 GND! VDD! _GENERATED_1440 _GENERATED_1439 261 279 sram_filler $T=9350 4620 0 0 $X=9354 $Y=4620
XX30BB92C5482 GND! VDD! _GENERATED_1442 _GENERATED_1441 263 VDD! sram_filler $T=9350 5544 0 0 $X=9354 $Y=5544
XX30BB92C5483 GND! VDD! _GENERATED_1444 _GENERATED_1443 264 VDD! sram_filler $T=9350 6468 0 0 $X=9354 $Y=6468
XX30BB92C5484 GND! VDD! GND! _GENERATED_1445 267 283 sram_filler $T=9350 11088 0 0 $X=9354 $Y=11088
XX30BB92C5485 GND! VDD! GND! _GENERATED_1446 268 287 sram_filler $T=9350 12012 0 0 $X=9354 $Y=12012
XX30BB92C5486 GND! VDD! GND! _GENERATED_1447 270 285 sram_filler $T=9350 13860 0 0 $X=9354 $Y=13860
XX30BB92C5487 GND! VDD! GND! _GENERATED_1448 269 286 sram_filler $T=9350 12936 0 0 $X=9354 $Y=12936
XX30BB92C5488 GND! VDD! GND! _GENERATED_1449 265 282 sram_filler $T=9350 9240 0 0 $X=9354 $Y=9240
XX30BB92C5489 GND! VDD! GND! _GENERATED_1450 266 284 sram_filler $T=9350 10164 0 0 $X=9354 $Y=10164
XX30BB92C5490 GND! VDD! GND! _GENERATED_1451 272 280 sram_filler $T=9350 8316 0 0 $X=9354 $Y=8316
XX30BB92C5491 GND! VDD! GND! _GENERATED_1452 262 281 sram_filler $T=9350 7392 0 0 $X=9354 $Y=7392
XX30BB92C5492 GND! VDD! GND! _GENERATED_1453 267 283 sram_filler $T=12374 11088 0 0 $X=12378 $Y=11088
XX30BB92C5493 GND! VDD! GND! _GENERATED_1454 268 287 sram_filler $T=12374 12012 0 0 $X=12378 $Y=12012
XX30BB92C5494 GND! VDD! GND! _GENERATED_1455 270 285 sram_filler $T=12374 13860 0 0 $X=12378 $Y=13860
XX30BB92C5495 GND! VDD! GND! _GENERATED_1456 269 286 sram_filler $T=12374 12936 0 0 $X=12378 $Y=12936
XX30BB92C5496 GND! VDD! GND! _GENERATED_1457 265 282 sram_filler $T=12374 9240 0 0 $X=12378 $Y=9240
XX30BB92C5497 GND! VDD! GND! _GENERATED_1458 266 284 sram_filler $T=12374 10164 0 0 $X=12378 $Y=10164
XX30BB92C5498 GND! VDD! GND! _GENERATED_1459 272 280 sram_filler $T=12374 8316 0 0 $X=12378 $Y=8316
XX30BB92C5499 GND! VDD! GND! _GENERATED_1460 262 281 sram_filler $T=12374 7392 0 0 $X=12378 $Y=7392
XX30BB92C5500 GND! VDD! GND! _GENERATED_1461 262 281 sram_filler $T=18422 7392 0 0 $X=18426 $Y=7392
XX30BB92C5501 GND! VDD! GND! _GENERATED_1462 272 280 sram_filler $T=18422 8316 0 0 $X=18426 $Y=8316
XX30BB92C5502 GND! VDD! GND! _GENERATED_1463 266 284 sram_filler $T=18422 10164 0 0 $X=18426 $Y=10164
XX30BB92C5503 GND! VDD! GND! _GENERATED_1464 265 282 sram_filler $T=18422 9240 0 0 $X=18426 $Y=9240
XX30BB92C5504 GND! VDD! GND! _GENERATED_1465 269 286 sram_filler $T=18422 12936 0 0 $X=18426 $Y=12936
XX30BB92C5505 GND! VDD! GND! _GENERATED_1466 270 285 sram_filler $T=18422 13860 0 0 $X=18426 $Y=13860
XX30BB92C5506 GND! VDD! GND! _GENERATED_1467 268 287 sram_filler $T=18422 12012 0 0 $X=18426 $Y=12012
XX30BB92C5507 GND! VDD! GND! _GENERATED_1468 267 283 sram_filler $T=18422 11088 0 0 $X=18426 $Y=11088
XX30BB92C5508 GND! VDD! GND! _GENERATED_1469 267 283 sram_filler $T=15398 11088 0 0 $X=15402 $Y=11088
XX30BB92C5509 GND! VDD! GND! _GENERATED_1470 268 287 sram_filler $T=15398 12012 0 0 $X=15402 $Y=12012
XX30BB92C5510 GND! VDD! GND! _GENERATED_1471 270 285 sram_filler $T=15398 13860 0 0 $X=15402 $Y=13860
XX30BB92C5511 GND! VDD! GND! _GENERATED_1472 269 286 sram_filler $T=15398 12936 0 0 $X=15402 $Y=12936
XX30BB92C5512 GND! VDD! GND! _GENERATED_1473 265 282 sram_filler $T=15398 9240 0 0 $X=15402 $Y=9240
XX30BB92C5513 GND! VDD! GND! _GENERATED_1474 266 284 sram_filler $T=15398 10164 0 0 $X=15402 $Y=10164
XX30BB92C5514 GND! VDD! GND! _GENERATED_1475 272 280 sram_filler $T=15398 8316 0 0 $X=15402 $Y=8316
XX30BB92C5515 GND! VDD! GND! _GENERATED_1476 262 281 sram_filler $T=15398 7392 0 0 $X=15402 $Y=7392
XX30BB92C5516 GND! VDD! _GENERATED_1478 _GENERATED_1477 257 276 sram_filler $T=6778 1050 0 180 $X=6330 $Y=460
XX30BB92C5517 GND! VDD! _GENERATED_1479 GND! 257 276 sram_filler $T=6442 1050 0 180 $X=5994 $Y=460
XX30BB92C5518 GND! VDD! VDD! _GENERATED_1480 257 276 sram_filler $T=6274 1050 0 180 $X=5826 $Y=460
XX30BB92C5519 GND! VDD! _GENERATED_1482 _GENERATED_1481 257 276 sram_filler $T=5938 1050 0 180 $X=5489 $Y=460
XX30BB92C5520 GND! VDD! _GENERATED_1484 _GENERATED_1483 257 276 sram_filler $T=394 1050 0 180 $X=-53 $Y=460
XX30BB92C5521 GND! VDD! _GENERATED_1486 _GENERATED_1485 257 276 sram_filler $T=730 1050 0 180 $X=282 $Y=460
XX30BB92C5522 GND! VDD! _GENERATED_1488 _GENERATED_1487 257 276 sram_filler $T=1402 1050 0 180 $X=954 $Y=460
XX30BB92C5523 GND! VDD! _GENERATED_1490 _GENERATED_1489 257 276 sram_filler $T=1066 1050 0 180 $X=618 $Y=460
XX30BB92C5524 GND! VDD! _GENERATED_1492 _GENERATED_1491 259 277 sram_filler $T=394 1974 0 180 $X=-53 $Y=1384
XX30BB92C5525 GND! VDD! _GENERATED_1494 _GENERATED_1493 259 277 sram_filler $T=730 1974 0 180 $X=282 $Y=1384
XX30BB92C5526 GND! VDD! _GENERATED_1496 _GENERATED_1495 259 277 sram_filler $T=1402 1974 0 180 $X=954 $Y=1384
XX30BB92C5527 GND! VDD! _GENERATED_1498 _GENERATED_1497 259 277 sram_filler $T=1066 1974 0 180 $X=618 $Y=1384
XX30BB92C5528 GND! VDD! _GENERATED_1500 _GENERATED_1499 258 278 sram_filler $T=1066 2898 0 180 $X=618 $Y=2308
XX30BB92C5529 GND! VDD! _GENERATED_1502 _GENERATED_1501 258 278 sram_filler $T=1402 2898 0 180 $X=954 $Y=2308
XX30BB92C5530 GND! VDD! _GENERATED_1504 _GENERATED_1503 258 278 sram_filler $T=730 2898 0 180 $X=282 $Y=2308
XX30BB92C5531 GND! VDD! _GENERATED_1506 _GENERATED_1505 258 278 sram_filler $T=394 2898 0 180 $X=-53 $Y=2308
XX30BB92C5532 GND! VDD! _GENERATED_1508 _GENERATED_1507 260 275 sram_filler $T=1066 3822 0 180 $X=618 $Y=3232
XX30BB92C5533 GND! VDD! _GENERATED_1510 _GENERATED_1509 260 275 sram_filler $T=1402 3822 0 180 $X=954 $Y=3232
XX30BB92C5534 GND! VDD! _GENERATED_1512 _GENERATED_1511 260 275 sram_filler $T=730 3822 0 180 $X=282 $Y=3232
XX30BB92C5535 GND! VDD! _GENERATED_1514 _GENERATED_1513 260 275 sram_filler $T=394 3822 0 180 $X=-53 $Y=3232
XX30BB92C5536 GND! VDD! _GENERATED_1516 _GENERATED_1515 258 278 sram_filler $T=18034 2898 0 180 $X=17586 $Y=2308
XX30BB92C5537 GND! VDD! _GENERATED_1518 _GENERATED_1517 258 278 sram_filler $T=18370 2898 0 180 $X=17922 $Y=2308
XX30BB92C5538 GND! VDD! 28 _GENERATED_1519 258 278 sram_filler $T=18706 2898 0 180 $X=18258 $Y=2308
XX30BB92C5539 GND! VDD! _GENERATED_1521 _GENERATED_1520 258 278 sram_filler $T=16690 2898 0 180 $X=16242 $Y=2308
XX30BB92C5540 GND! VDD! _GENERATED_1523 _GENERATED_1522 258 278 sram_filler $T=17026 2898 0 180 $X=16578 $Y=2308
XX30BB92C5541 GND! VDD! _GENERATED_1525 _GENERATED_1524 258 278 sram_filler $T=17362 2898 0 180 $X=16914 $Y=2308
XX30BB92C5542 GND! VDD! _GENERATED_1527 _GENERATED_1526 258 278 sram_filler $T=17698 2898 0 180 $X=17250 $Y=2308
XX30BB92C5543 GND! VDD! VDD! _GENERATED_1528 259 277 sram_filler $T=6610 1974 0 180 $X=6162 $Y=1384
XX30BB92C5544 GND! VDD! _GENERATED_1530 _GENERATED_1529 259 277 sram_filler $T=6274 1974 0 180 $X=5826 $Y=1384
XX30BB92C5545 GND! VDD! _GENERATED_1532 _GENERATED_1531 259 277 sram_filler $T=5938 1974 0 180 $X=5489 $Y=1384
XX30BB92C5546 GND! VDD! _GENERATED_1533 GND! 259 277 sram_filler $T=6778 1974 0 180 $X=6330 $Y=1384
XX30BB92C5547 GND! VDD! _GENERATED_1535 _GENERATED_1534 258 278 sram_filler $T=11986 2898 0 180 $X=11538 $Y=2308
XX30BB92C5548 GND! VDD! _GENERATED_1537 _GENERATED_1536 258 278 sram_filler $T=12322 2898 0 180 $X=11874 $Y=2308
XX30BB92C5549 GND! VDD! _GENERATED_1539 _GENERATED_1538 258 278 sram_filler $T=12658 2898 0 180 $X=12209 $Y=2308
XX30BB92C5550 GND! VDD! _GENERATED_1541 _GENERATED_1540 258 278 sram_filler $T=12994 2898 0 180 $X=12546 $Y=2308
XX30BB92C5551 GND! VDD! _GENERATED_1543 _GENERATED_1542 258 278 sram_filler $T=13330 2898 0 180 $X=12882 $Y=2308
XX30BB92C5552 GND! VDD! _GENERATED_1545 _GENERATED_1544 258 278 sram_filler $T=11314 2898 0 180 $X=10866 $Y=2308
XX30BB92C5553 GND! VDD! _GENERATED_1547 _GENERATED_1546 258 278 sram_filler $T=11650 2898 0 180 $X=11202 $Y=2308
XX30BB92C5554 GND! VDD! _GENERATED_1549 _GENERATED_1548 258 278 sram_filler $T=13666 2898 0 180 $X=13218 $Y=2308
XX30BB92C5555 GND! VDD! _GENERATED_1551 _GENERATED_1550 258 278 sram_filler $T=14002 2898 0 180 $X=13554 $Y=2308
XX30BB92C5556 GND! VDD! _GENERATED_1553 _GENERATED_1552 258 278 sram_filler $T=14338 2898 0 180 $X=13890 $Y=2308
XX30BB92C5557 GND! VDD! _GENERATED_1555 _GENERATED_1554 258 278 sram_filler $T=14674 2898 0 180 $X=14226 $Y=2308
XX30BB92C5558 GND! VDD! _GENERATED_1557 _GENERATED_1556 258 278 sram_filler $T=15010 2898 0 180 $X=14562 $Y=2308
XX30BB92C5559 GND! VDD! _GENERATED_1559 _GENERATED_1558 258 278 sram_filler $T=15346 2898 0 180 $X=14898 $Y=2308
XX30BB92C5560 GND! VDD! _GENERATED_1561 _GENERATED_1560 258 278 sram_filler $T=16018 2898 0 180 $X=15570 $Y=2308
XX30BB92C5561 GND! VDD! _GENERATED_1563 _GENERATED_1562 258 278 sram_filler $T=15682 2898 0 180 $X=15234 $Y=2308
XX30BB92C5562 GND! VDD! _GENERATED_1565 _GENERATED_1564 258 278 sram_filler $T=16354 2898 0 180 $X=15905 $Y=2308
XX30BB92C5563 GND! VDD! _GENERATED_1567 _GENERATED_1566 258 278 sram_filler $T=9970 2898 0 180 $X=9522 $Y=2308
XX30BB92C5564 GND! VDD! _GENERATED_1569 _GENERATED_1568 258 278 sram_filler $T=10306 2898 0 180 $X=9858 $Y=2308
XX30BB92C5565 GND! VDD! _GENERATED_1571 _GENERATED_1570 258 278 sram_filler $T=10642 2898 0 180 $X=10193 $Y=2308
XX30BB92C5566 GND! VDD! _GENERATED_1573 _GENERATED_1572 258 278 sram_filler $T=10978 2898 0 180 $X=10530 $Y=2308
XX30BB92C5567 GND! VDD! _GENERATED_1575 _GENERATED_1574 258 278 sram_filler $T=9634 2898 0 180 $X=9186 $Y=2308
XX30BB92C5568 GND! VDD! _GENERATED_1577 _GENERATED_1576 258 278 sram_filler $T=9298 2898 0 180 $X=8850 $Y=2308
XX30BB92C5569 GND! VDD! _GENERATED_1579 _GENERATED_1578 258 278 sram_filler $T=8962 2898 0 180 $X=8514 $Y=2308
XX30BB92C5570 GND! VDD! _GENERATED_1581 _GENERATED_1580 258 278 sram_filler $T=8626 2898 0 180 $X=8177 $Y=2308
XX30BB92C5571 GND! VDD! _GENERATED_1583 _GENERATED_1582 258 278 sram_filler $T=6946 2898 0 180 $X=6497 $Y=2308
XX30BB92C5572 GND! VDD! _GENERATED_1585 _GENERATED_1584 258 278 sram_filler $T=6610 2898 0 180 $X=6162 $Y=2308
XX30BB92C5573 GND! VDD! _GENERATED_1587 _GENERATED_1586 258 278 sram_filler $T=6274 2898 0 180 $X=5826 $Y=2308
XX30BB92C5574 GND! VDD! _GENERATED_1589 _GENERATED_1588 258 278 sram_filler $T=5938 2898 0 180 $X=5489 $Y=2308
XX30BB92C5575 GND! VDD! _GENERATED_1591 _GENERATED_1590 258 278 sram_filler $T=8290 2898 0 180 $X=7842 $Y=2308
XX30BB92C5576 GND! VDD! _GENERATED_1593 _GENERATED_1592 258 278 sram_filler $T=7954 2898 0 180 $X=7505 $Y=2308
XX30BB92C5577 GND! VDD! _GENERATED_1595 _GENERATED_1594 258 278 sram_filler $T=7618 2898 0 180 $X=7170 $Y=2308
XX30BB92C5578 GND! VDD! _GENERATED_1597 _GENERATED_1596 258 278 sram_filler $T=7282 2898 0 180 $X=6834 $Y=2308
XX30BB92C5579 GND! VDD! _GENERATED_1599 _GENERATED_1598 264 VDD! sram_filler $T=15850 6594 0 180 $X=15402 $Y=6004
XX30BB92C5580 GND! VDD! _GENERATED_1601 _GENERATED_1600 263 279 sram_filler $T=15850 5670 0 180 $X=15402 $Y=5080
XX30BB92C5581 GND! VDD! _GENERATED_1603 _GENERATED_1602 261 274 sram_filler $T=15850 4746 0 180 $X=15402 $Y=4156
XX30BB92C5582 GND! VDD! _GENERATED_1605 _GENERATED_1604 260 275 sram_filler $T=15850 3822 0 180 $X=15402 $Y=3232
XX30BB92C5583 GND! VDD! _GENERATED_1607 _GENERATED_1606 261 274 sram_filler $T=12826 4746 0 180 $X=12378 $Y=4156
XX30BB92C5584 GND! VDD! _GENERATED_1609 _GENERATED_1608 260 275 sram_filler $T=12826 3822 0 180 $X=12378 $Y=3232
XX30BB92C5585 GND! VDD! _GENERATED_1611 _GENERATED_1610 263 279 sram_filler $T=12826 5670 0 180 $X=12378 $Y=5080
XX30BB92C5586 GND! VDD! _GENERATED_1613 _GENERATED_1612 264 VDD! sram_filler $T=12826 6594 0 180 $X=12378 $Y=6004
XX30BB92C5587 GND! VDD! _GENERATED_1615 _GENERATED_1614 260 275 sram_filler $T=9802 3822 0 180 $X=9354 $Y=3232
XX30BB92C5588 GND! VDD! _GENERATED_1617 _GENERATED_1616 261 274 sram_filler $T=9802 4746 0 180 $X=9354 $Y=4156
XX30BB92C5589 GND! VDD! _GENERATED_1619 _GENERATED_1618 263 279 sram_filler $T=9802 5670 0 180 $X=9354 $Y=5080
XX30BB92C5590 GND! VDD! _GENERATED_1621 _GENERATED_1620 264 VDD! sram_filler $T=9802 6594 0 180 $X=9354 $Y=6004
XX30BB92C5591 GND! VDD! VDD! _GENERATED_1622 262 VDD! sram_filler $T=5938 7518 0 180 $X=5489 $Y=6928
XX30BB92C5592 GND! VDD! _GENERATED_1623 GND! 262 VDD! sram_filler $T=6106 7518 0 180 $X=5657 $Y=6928
XX30BB92C5593 GND! VDD! _GENERATED_1625 _GENERATED_1624 262 VDD! sram_filler $T=6442 7518 0 180 $X=5994 $Y=6928
XX30BB92C5594 GND! VDD! VDD! _GENERATED_1626 261 274 sram_filler $T=394 4746 0 180 $X=-53 $Y=4156
XX30BB92C5595 GND! VDD! _GENERATED_1628 _GENERATED_1627 261 274 sram_filler $T=2914 4746 0 180 $X=2466 $Y=4156
XX30BB92C5596 GND! VDD! _GENERATED_1630 _GENERATED_1629 261 274 sram_filler $T=2578 4746 0 180 $X=2130 $Y=4156
XX30BB92C5597 GND! VDD! _GENERATED_1632 _GENERATED_1631 261 274 sram_filler $T=1906 4746 0 180 $X=1458 $Y=4156
XX30BB92C5598 GND! VDD! _GENERATED_1634 _GENERATED_1633 261 274 sram_filler $T=2242 4746 0 180 $X=1794 $Y=4156
XX30BB92C5599 GND! VDD! _GENERATED_1636 _GENERATED_1635 261 274 sram_filler $T=1234 4746 0 180 $X=786 $Y=4156
XX30BB92C5600 GND! VDD! _GENERATED_1638 _GENERATED_1637 261 274 sram_filler $T=1570 4746 0 180 $X=1122 $Y=4156
XX30BB92C5601 GND! VDD! _GENERATED_1639 GND! 261 274 sram_filler $T=562 4746 0 180 $X=114 $Y=4156
XX30BB92C5602 GND! VDD! _GENERATED_1641 _GENERATED_1640 261 274 sram_filler $T=898 4746 0 180 $X=450 $Y=4156
XX30BB92C5603 GND! VDD! _GENERATED_1643 _GENERATED_1642 261 274 sram_filler $T=3586 4746 0 180 $X=3138 $Y=4156
XX30BB92C5604 GND! VDD! _GENERATED_1645 _GENERATED_1644 261 274 sram_filler $T=3250 4746 0 180 $X=2802 $Y=4156
XX30BB92C5605 GND! VDD! _GENERATED_1647 _GENERATED_1646 261 274 sram_filler $T=4258 4746 0 180 $X=3810 $Y=4156
XX30BB92C5606 GND! VDD! _GENERATED_1649 _GENERATED_1648 261 274 sram_filler $T=3922 4746 0 180 $X=3474 $Y=4156
XX30BB92C5607 GND! VDD! _GENERATED_1651 _GENERATED_1650 261 274 sram_filler $T=4930 4746 0 180 $X=4481 $Y=4156
XX30BB92C5608 GND! VDD! _GENERATED_1653 _GENERATED_1652 261 274 sram_filler $T=4594 4746 0 180 $X=4146 $Y=4156
XX30BB92C5609 GND! VDD! _GENERATED_1655 _GENERATED_1654 261 274 sram_filler $T=5266 4746 0 180 $X=4818 $Y=4156
XX30BB92C5610 GND! VDD! _GENERATED_1657 _GENERATED_1656 261 274 sram_filler $T=5602 4746 0 180 $X=5154 $Y=4156
XX30BB92C5611 GND! VDD! _GENERATED_1659 _GENERATED_1658 262 VDD! sram_filler $T=6778 7518 0 180 $X=6330 $Y=6928
XX30BB92C5612 GND! VDD! GND! _GENERATED_1660 268 283 sram_filler $T=9350 12138 1 0 $X=9354 $Y=11548
XX30BB92C5613 GND! VDD! GND! _GENERATED_1661 269 287 sram_filler $T=9350 13062 1 0 $X=9354 $Y=12472
XX30BB92C5614 GND! VDD! GND! _GENERATED_1662 271 285 sram_filler $T=9350 14910 1 0 $X=9354 $Y=14320
XX30BB92C5615 GND! VDD! GND! _GENERATED_1663 270 286 sram_filler $T=9350 13986 1 0 $X=9354 $Y=13396
XX30BB92C5616 GND! VDD! GND! _GENERATED_1664 266 282 sram_filler $T=9350 10290 1 0 $X=9354 $Y=9700
XX30BB92C5617 GND! VDD! GND! _GENERATED_1665 267 284 sram_filler $T=9350 11214 1 0 $X=9354 $Y=10624
XX30BB92C5618 GND! VDD! GND! _GENERATED_1666 265 280 sram_filler $T=9350 9366 1 0 $X=9354 $Y=8776
XX30BB92C5619 GND! VDD! GND! _GENERATED_1667 272 281 sram_filler $T=9350 8442 1 0 $X=9354 $Y=7852
XX30BB92C5620 GND! VDD! GND! _GENERATED_1668 268 283 sram_filler $T=12374 12138 1 0 $X=12378 $Y=11548
XX30BB92C5621 GND! VDD! GND! _GENERATED_1669 269 287 sram_filler $T=12374 13062 1 0 $X=12378 $Y=12472
XX30BB92C5622 GND! VDD! GND! _GENERATED_1670 271 285 sram_filler $T=12374 14910 1 0 $X=12378 $Y=14320
XX30BB92C5623 GND! VDD! GND! _GENERATED_1671 270 286 sram_filler $T=12374 13986 1 0 $X=12378 $Y=13396
XX30BB92C5624 GND! VDD! GND! _GENERATED_1672 266 282 sram_filler $T=12374 10290 1 0 $X=12378 $Y=9700
XX30BB92C5625 GND! VDD! GND! _GENERATED_1673 267 284 sram_filler $T=12374 11214 1 0 $X=12378 $Y=10624
XX30BB92C5626 GND! VDD! GND! _GENERATED_1674 265 280 sram_filler $T=12374 9366 1 0 $X=12378 $Y=8776
XX30BB92C5627 GND! VDD! GND! _GENERATED_1675 272 281 sram_filler $T=12374 8442 1 0 $X=12378 $Y=7852
XX30BB92C5628 GND! VDD! GND! _GENERATED_1676 272 281 sram_filler $T=18422 8442 1 0 $X=18426 $Y=7852
XX30BB92C5629 GND! VDD! GND! _GENERATED_1677 265 280 sram_filler $T=18422 9366 1 0 $X=18426 $Y=8776
XX30BB92C5630 GND! VDD! GND! _GENERATED_1678 267 284 sram_filler $T=18422 11214 1 0 $X=18426 $Y=10624
XX30BB92C5631 GND! VDD! GND! _GENERATED_1679 266 282 sram_filler $T=18422 10290 1 0 $X=18426 $Y=9700
XX30BB92C5632 GND! VDD! GND! _GENERATED_1680 270 286 sram_filler $T=18422 13986 1 0 $X=18426 $Y=13396
XX30BB92C5633 GND! VDD! GND! _GENERATED_1681 271 285 sram_filler $T=18422 14910 1 0 $X=18426 $Y=14320
XX30BB92C5634 GND! VDD! GND! _GENERATED_1682 269 287 sram_filler $T=18422 13062 1 0 $X=18426 $Y=12472
XX30BB92C5635 GND! VDD! GND! _GENERATED_1683 268 283 sram_filler $T=18422 12138 1 0 $X=18426 $Y=11548
XX30BB92C5636 GND! VDD! GND! _GENERATED_1684 268 283 sram_filler $T=15398 12138 1 0 $X=15402 $Y=11548
XX30BB92C5637 GND! VDD! GND! _GENERATED_1685 269 287 sram_filler $T=15398 13062 1 0 $X=15402 $Y=12472
XX30BB92C5638 GND! VDD! GND! _GENERATED_1686 271 285 sram_filler $T=15398 14910 1 0 $X=15402 $Y=14320
XX30BB92C5639 GND! VDD! GND! _GENERATED_1687 270 286 sram_filler $T=15398 13986 1 0 $X=15402 $Y=13396
XX30BB92C5640 GND! VDD! GND! _GENERATED_1688 266 282 sram_filler $T=15398 10290 1 0 $X=15402 $Y=9700
XX30BB92C5641 GND! VDD! GND! _GENERATED_1689 267 284 sram_filler $T=15398 11214 1 0 $X=15402 $Y=10624
XX30BB92C5642 GND! VDD! GND! _GENERATED_1690 265 280 sram_filler $T=15398 9366 1 0 $X=15402 $Y=8776
XX30BB92C5643 GND! VDD! GND! _GENERATED_1691 272 281 sram_filler $T=15398 8442 1 0 $X=15402 $Y=7852
XX30BB92C5644 GND! VDD! GND! 9 373 140 12 103 177 104 265 
+	266 282 sram_6t $T=6690 9240 0 0 $X=6666 $Y=9240
XX30BB92C5645 GND! VDD! GND! 9 341 487 8 98 133 99 262 
+	272 281 sram_6t $T=8706 7392 0 0 $X=8682 $Y=7392
XX30BB92C5646 GND! VDD! GND! 9 342 488 10 98 134 99 262 
+	272 281 sram_6t $T=8034 7392 0 0 $X=8010 $Y=7392
XX30BB92C5647 GND! VDD! GND! 9 343 489 11 98 135 99 262 
+	272 281 sram_6t $T=7362 7392 0 0 $X=7338 $Y=7392
XX30BB92C5648 GND! VDD! GND! 9 344 135 11 99 136 103 272 
+	265 280 sram_6t $T=7362 8316 0 0 $X=7338 $Y=8316
XX30BB92C5649 GND! VDD! GND! 9 345 134 10 99 137 103 272 
+	265 280 sram_6t $T=8034 8316 0 0 $X=8010 $Y=8316
XX30BB92C5650 GND! VDD! GND! 9 346 133 8 99 138 103 272 
+	265 280 sram_6t $T=8706 8316 0 0 $X=8682 $Y=8316
XX30BB92C5651 GND! VDD! GND! 9 347 490 12 98 139 99 262 
+	272 281 sram_6t $T=6690 7392 0 0 $X=6666 $Y=7392
XX30BB92C5652 GND! VDD! GND! 9 348 139 12 99 140 103 272 
+	265 280 sram_6t $T=6690 8316 0 0 $X=6666 $Y=8316
XX30BB92C5653 GND! VDD! GND! 9 374 136 11 103 178 104 265 
+	266 282 sram_6t $T=7362 9240 0 0 $X=7338 $Y=9240
XX30BB92C5654 GND! VDD! GND! 9 375 137 10 103 179 104 265 
+	266 282 sram_6t $T=8034 9240 0 0 $X=8010 $Y=9240
XX30BB92C5655 GND! VDD! GND! 9 376 138 8 103 180 104 265 
+	266 282 sram_6t $T=8706 9240 0 0 $X=8682 $Y=9240
XX30BB92C5656 GND! VDD! GND! 9 377 177 12 104 181 105 266 
+	267 284 sram_6t $T=6690 10164 0 0 $X=6666 $Y=10164
XX30BB92C5657 GND! VDD! GND! 9 378 180 8 104 182 105 266 
+	267 284 sram_6t $T=8706 10164 0 0 $X=8682 $Y=10164
XX30BB92C5658 GND! VDD! GND! 9 379 179 10 104 183 105 266 
+	267 284 sram_6t $T=8034 10164 0 0 $X=8010 $Y=10164
XX30BB92C5659 GND! VDD! GND! 9 380 178 11 104 184 105 266 
+	267 284 sram_6t $T=7362 10164 0 0 $X=7338 $Y=10164
XX30BB92C5660 GND! VDD! GND! 9 381 182 8 105 185 106 267 
+	268 283 sram_6t $T=8706 11088 0 0 $X=8682 $Y=11088
XX30BB92C5661 GND! VDD! GND! 9 382 183 10 105 186 106 267 
+	268 283 sram_6t $T=8034 11088 0 0 $X=8010 $Y=11088
XX30BB92C5662 GND! VDD! GND! 9 383 184 11 105 187 106 267 
+	268 283 sram_6t $T=7362 11088 0 0 $X=7338 $Y=11088
XX30BB92C5663 GND! VDD! GND! 9 384 181 12 105 188 106 267 
+	268 283 sram_6t $T=6690 11088 0 0 $X=6666 $Y=11088
XX30BB92C5664 GND! VDD! GND! 9 421 187 11 106 189 107 268 
+	269 287 sram_6t $T=7362 12012 0 0 $X=7338 $Y=12012
XX30BB92C5665 GND! VDD! GND! 9 422 186 10 106 190 107 268 
+	269 287 sram_6t $T=8034 12012 0 0 $X=8010 $Y=12012
XX30BB92C5666 GND! VDD! GND! 9 423 185 8 106 191 107 268 
+	269 287 sram_6t $T=8706 12012 0 0 $X=8682 $Y=12012
XX30BB92C5667 GND! VDD! GND! 9 424 188 12 106 192 107 268 
+	269 287 sram_6t $T=6690 12012 0 0 $X=6666 $Y=12012
XX30BB92C5668 GND! VDD! GND! 9 425 192 12 107 193 108 269 
+	270 286 sram_6t $T=6690 12936 0 0 $X=6666 $Y=12936
XX30BB92C5669 GND! VDD! GND! 9 426 189 11 107 194 108 269 
+	270 286 sram_6t $T=7362 12936 0 0 $X=7338 $Y=12936
XX30BB92C5670 GND! VDD! GND! 9 427 190 10 107 195 108 269 
+	270 286 sram_6t $T=8034 12936 0 0 $X=8010 $Y=12936
XX30BB92C5671 GND! VDD! GND! 9 428 191 8 107 196 108 269 
+	270 286 sram_6t $T=8706 12936 0 0 $X=8682 $Y=12936
XX30BB92C5672 GND! VDD! GND! 9 429 193 12 108 512 513 270 
+	271 285 sram_6t $T=6690 13860 0 0 $X=6666 $Y=13860
XX30BB92C5673 GND! VDD! GND! 9 430 196 8 108 518 519 270 
+	271 285 sram_6t $T=8706 13860 0 0 $X=8682 $Y=13860
XX30BB92C5674 GND! VDD! GND! 9 431 195 10 108 516 517 270 
+	271 285 sram_6t $T=8034 13860 0 0 $X=8010 $Y=13860
XX30BB92C5675 GND! VDD! GND! 9 432 194 11 108 514 515 270 
+	271 285 sram_6t $T=7362 13860 0 0 $X=7338 $Y=13860
XX30BB92C5676 GND! VDD! GND! 14 433 197 15 108 522 523 270 
+	271 285 sram_6t $T=10386 13860 0 0 $X=10362 $Y=13860
XX30BB92C5677 GND! VDD! GND! 14 434 198 16 108 524 525 270 
+	271 285 sram_6t $T=11058 13860 0 0 $X=11034 $Y=13860
XX30BB92C5678 GND! VDD! GND! 14 435 199 17 108 526 527 270 
+	271 285 sram_6t $T=11730 13860 0 0 $X=11706 $Y=13860
XX30BB92C5679 GND! VDD! GND! 14 436 200 13 108 520 521 270 
+	271 285 sram_6t $T=9714 13860 0 0 $X=9690 $Y=13860
XX30BB92C5680 GND! VDD! GND! 14 437 201 17 107 199 108 269 
+	270 286 sram_6t $T=11730 12936 0 0 $X=11706 $Y=12936
XX30BB92C5681 GND! VDD! GND! 14 438 202 16 107 198 108 269 
+	270 286 sram_6t $T=11058 12936 0 0 $X=11034 $Y=12936
XX30BB92C5682 GND! VDD! GND! 14 439 203 15 107 197 108 269 
+	270 286 sram_6t $T=10386 12936 0 0 $X=10362 $Y=12936
XX30BB92C5683 GND! VDD! GND! 14 440 204 13 107 200 108 269 
+	270 286 sram_6t $T=9714 12936 0 0 $X=9690 $Y=12936
XX30BB92C5684 GND! VDD! GND! 14 441 205 13 106 204 107 268 
+	269 287 sram_6t $T=9714 12012 0 0 $X=9690 $Y=12012
XX30BB92C5685 GND! VDD! GND! 14 442 206 17 106 201 107 268 
+	269 287 sram_6t $T=11730 12012 0 0 $X=11706 $Y=12012
XX30BB92C5686 GND! VDD! GND! 14 443 207 16 106 202 107 268 
+	269 287 sram_6t $T=11058 12012 0 0 $X=11034 $Y=12012
XX30BB92C5687 GND! VDD! GND! 14 444 208 15 106 203 107 268 
+	269 287 sram_6t $T=10386 12012 0 0 $X=10362 $Y=12012
XX30BB92C5688 GND! VDD! GND! 14 385 209 13 105 205 106 267 
+	268 283 sram_6t $T=9714 11088 0 0 $X=9690 $Y=11088
XX30BB92C5689 GND! VDD! GND! 14 386 210 15 105 208 106 267 
+	268 283 sram_6t $T=10386 11088 0 0 $X=10362 $Y=11088
XX30BB92C5690 GND! VDD! GND! 14 387 211 16 105 207 106 267 
+	268 283 sram_6t $T=11058 11088 0 0 $X=11034 $Y=11088
XX30BB92C5691 GND! VDD! GND! 14 388 212 17 105 206 106 267 
+	268 283 sram_6t $T=11730 11088 0 0 $X=11706 $Y=11088
XX30BB92C5692 GND! VDD! GND! 14 389 213 15 104 210 105 266 
+	267 284 sram_6t $T=10386 10164 0 0 $X=10362 $Y=10164
XX30BB92C5693 GND! VDD! GND! 14 390 214 16 104 211 105 266 
+	267 284 sram_6t $T=11058 10164 0 0 $X=11034 $Y=10164
XX30BB92C5694 GND! VDD! GND! 14 391 215 17 104 212 105 266 
+	267 284 sram_6t $T=11730 10164 0 0 $X=11706 $Y=10164
XX30BB92C5695 GND! VDD! GND! 14 392 216 13 104 209 105 266 
+	267 284 sram_6t $T=9714 10164 0 0 $X=9690 $Y=10164
XX30BB92C5696 GND! VDD! GND! 14 393 152 17 103 215 104 265 
+	266 282 sram_6t $T=11730 9240 0 0 $X=11706 $Y=9240
XX30BB92C5697 GND! VDD! GND! 14 394 150 16 103 214 104 265 
+	266 282 sram_6t $T=11058 9240 0 0 $X=11034 $Y=9240
XX30BB92C5698 GND! VDD! GND! 14 395 148 15 103 213 104 265 
+	266 282 sram_6t $T=10386 9240 0 0 $X=10362 $Y=9240
XX30BB92C5699 GND! VDD! GND! 14 396 146 13 103 216 104 265 
+	266 282 sram_6t $T=9714 9240 0 0 $X=9690 $Y=9240
XX30BB92C5700 GND! VDD! GND! 14 349 145 13 99 146 103 272 
+	265 280 sram_6t $T=9714 8316 0 0 $X=9690 $Y=8316
XX30BB92C5701 GND! VDD! GND! 14 350 147 15 99 148 103 272 
+	265 280 sram_6t $T=10386 8316 0 0 $X=10362 $Y=8316
XX30BB92C5702 GND! VDD! GND! 14 351 149 16 99 150 103 272 
+	265 280 sram_6t $T=11058 8316 0 0 $X=11034 $Y=8316
XX30BB92C5703 GND! VDD! GND! 14 352 151 17 99 152 103 272 
+	265 280 sram_6t $T=11730 8316 0 0 $X=11706 $Y=8316
XX30BB92C5704 GND! VDD! GND! 14 353 491 17 98 151 99 262 
+	272 281 sram_6t $T=11730 7392 0 0 $X=11706 $Y=7392
XX30BB92C5705 GND! VDD! GND! 14 354 492 16 98 149 99 262 
+	272 281 sram_6t $T=11058 7392 0 0 $X=11034 $Y=7392
XX30BB92C5706 GND! VDD! GND! 14 355 493 15 98 147 99 262 
+	272 281 sram_6t $T=10386 7392 0 0 $X=10362 $Y=7392
XX30BB92C5707 GND! VDD! GND! 14 356 494 13 98 145 99 262 
+	272 281 sram_6t $T=9714 7392 0 0 $X=9690 $Y=7392
XX30BB92C5708 GND! VDD! GND! 24 357 169 27 99 170 103 272 
+	265 280 sram_6t $T=17778 8316 0 0 $X=17753 $Y=8316
XX30BB92C5709 GND! VDD! GND! 24 358 171 26 99 172 103 272 
+	265 280 sram_6t $T=17106 8316 0 0 $X=17082 $Y=8316
XX30BB92C5710 GND! VDD! GND! 24 359 173 25 99 174 103 272 
+	265 280 sram_6t $T=16434 8316 0 0 $X=16410 $Y=8316
XX30BB92C5711 GND! VDD! GND! 24 360 175 23 99 176 103 272 
+	265 280 sram_6t $T=15762 8316 0 0 $X=15738 $Y=8316
XX30BB92C5712 GND! VDD! GND! 24 397 176 23 103 237 104 265 
+	266 282 sram_6t $T=15762 9240 0 0 $X=15738 $Y=9240
XX30BB92C5713 GND! VDD! GND! 24 398 174 25 103 238 104 265 
+	266 282 sram_6t $T=16434 9240 0 0 $X=16410 $Y=9240
XX30BB92C5714 GND! VDD! GND! 24 399 172 26 103 239 104 265 
+	266 282 sram_6t $T=17106 9240 0 0 $X=17082 $Y=9240
XX30BB92C5715 GND! VDD! GND! 24 400 170 27 103 240 104 265 
+	266 282 sram_6t $T=17778 9240 0 0 $X=17753 $Y=9240
XX30BB92C5716 GND! VDD! GND! 24 401 237 23 104 241 105 266 
+	267 284 sram_6t $T=15762 10164 0 0 $X=15738 $Y=10164
XX30BB92C5717 GND! VDD! GND! 24 402 240 27 104 242 105 266 
+	267 284 sram_6t $T=17778 10164 0 0 $X=17753 $Y=10164
XX30BB92C5718 GND! VDD! GND! 24 403 239 26 104 243 105 266 
+	267 284 sram_6t $T=17106 10164 0 0 $X=17082 $Y=10164
XX30BB92C5719 GND! VDD! GND! 24 404 238 25 104 244 105 266 
+	267 284 sram_6t $T=16434 10164 0 0 $X=16410 $Y=10164
XX30BB92C5720 GND! VDD! GND! 24 405 242 27 105 245 106 267 
+	268 283 sram_6t $T=17778 11088 0 0 $X=17753 $Y=11088
XX30BB92C5721 GND! VDD! GND! 24 406 243 26 105 246 106 267 
+	268 283 sram_6t $T=17106 11088 0 0 $X=17082 $Y=11088
XX30BB92C5722 GND! VDD! GND! 24 407 244 25 105 247 106 267 
+	268 283 sram_6t $T=16434 11088 0 0 $X=16410 $Y=11088
XX30BB92C5723 GND! VDD! GND! 24 408 241 23 105 248 106 267 
+	268 283 sram_6t $T=15762 11088 0 0 $X=15738 $Y=11088
XX30BB92C5724 GND! VDD! GND! 24 445 247 25 106 249 107 268 
+	269 287 sram_6t $T=16434 12012 0 0 $X=16410 $Y=12012
XX30BB92C5725 GND! VDD! GND! 24 446 246 26 106 250 107 268 
+	269 287 sram_6t $T=17106 12012 0 0 $X=17082 $Y=12012
XX30BB92C5726 GND! VDD! GND! 24 447 245 27 106 251 107 268 
+	269 287 sram_6t $T=17778 12012 0 0 $X=17753 $Y=12012
XX30BB92C5727 GND! VDD! GND! 24 448 248 23 106 252 107 268 
+	269 287 sram_6t $T=15762 12012 0 0 $X=15738 $Y=12012
XX30BB92C5728 GND! VDD! GND! 24 449 252 23 107 253 108 269 
+	270 286 sram_6t $T=15762 12936 0 0 $X=15738 $Y=12936
XX30BB92C5729 GND! VDD! GND! 24 450 249 25 107 254 108 269 
+	270 286 sram_6t $T=16434 12936 0 0 $X=16410 $Y=12936
XX30BB92C5730 GND! VDD! GND! 24 451 250 26 107 255 108 269 
+	270 286 sram_6t $T=17106 12936 0 0 $X=17082 $Y=12936
XX30BB92C5731 GND! VDD! GND! 24 452 251 27 107 256 108 269 
+	270 286 sram_6t $T=17778 12936 0 0 $X=17753 $Y=12936
XX30BB92C5732 GND! VDD! GND! 24 453 253 23 108 536 537 270 
+	271 285 sram_6t $T=15762 13860 0 0 $X=15738 $Y=13860
XX30BB92C5733 GND! VDD! GND! 24 454 256 27 108 542 543 270 
+	271 285 sram_6t $T=17778 13860 0 0 $X=17753 $Y=13860
XX30BB92C5734 GND! VDD! GND! 24 455 255 26 108 540 541 270 
+	271 285 sram_6t $T=17106 13860 0 0 $X=17082 $Y=13860
XX30BB92C5735 GND! VDD! GND! 24 456 254 25 108 538 539 270 
+	271 285 sram_6t $T=16434 13860 0 0 $X=16410 $Y=13860
XX30BB92C5736 GND! VDD! GND! 19 457 217 22 108 534 535 270 
+	271 285 sram_6t $T=14754 13860 0 0 $X=14730 $Y=13860
XX30BB92C5737 GND! VDD! GND! 19 458 218 22 107 217 108 269 
+	270 286 sram_6t $T=14754 12936 0 0 $X=14730 $Y=12936
XX30BB92C5738 GND! VDD! GND! 19 459 219 22 106 218 107 268 
+	269 287 sram_6t $T=14754 12012 0 0 $X=14730 $Y=12012
XX30BB92C5739 GND! VDD! GND! 19 409 220 22 105 219 106 267 
+	268 283 sram_6t $T=14754 11088 0 0 $X=14730 $Y=11088
XX30BB92C5740 GND! VDD! GND! 19 410 221 22 104 220 105 266 
+	267 284 sram_6t $T=14754 10164 0 0 $X=14730 $Y=10164
XX30BB92C5741 GND! VDD! GND! 19 411 158 22 103 221 104 265 
+	266 282 sram_6t $T=14754 9240 0 0 $X=14730 $Y=9240
XX30BB92C5742 GND! VDD! GND! 19 361 157 22 99 158 103 272 
+	265 280 sram_6t $T=14754 8316 0 0 $X=14730 $Y=8316
XX30BB92C5743 GND! VDD! GND! 24 362 497 23 98 175 99 262 
+	272 281 sram_6t $T=15762 7392 0 0 $X=15738 $Y=7392
XX30BB92C5744 GND! VDD! GND! 24 363 498 25 98 173 99 262 
+	272 281 sram_6t $T=16434 7392 0 0 $X=16410 $Y=7392
XX30BB92C5745 GND! VDD! GND! 24 364 499 26 98 171 99 262 
+	272 281 sram_6t $T=17106 7392 0 0 $X=17082 $Y=7392
XX30BB92C5746 GND! VDD! GND! 24 365 500 27 98 169 99 262 
+	272 281 sram_6t $T=17778 7392 0 0 $X=17753 $Y=7392
XX30BB92C5747 GND! VDD! GND! 19 460 222 20 108 530 531 270 
+	271 285 sram_6t $T=13410 13860 0 0 $X=13386 $Y=13860
XX30BB92C5748 GND! VDD! GND! 19 461 223 18 108 532 533 270 
+	271 285 sram_6t $T=14082 13860 0 0 $X=14058 $Y=13860
XX30BB92C5749 GND! VDD! GND! 19 462 224 21 108 528 529 270 
+	271 285 sram_6t $T=12738 13860 0 0 $X=12714 $Y=13860
XX30BB92C5750 GND! VDD! GND! 19 463 225 18 107 223 108 269 
+	270 286 sram_6t $T=14082 12936 0 0 $X=14058 $Y=12936
XX30BB92C5751 GND! VDD! GND! 19 464 226 20 107 222 108 269 
+	270 286 sram_6t $T=13410 12936 0 0 $X=13386 $Y=12936
XX30BB92C5752 GND! VDD! GND! 19 465 227 21 107 224 108 269 
+	270 286 sram_6t $T=12738 12936 0 0 $X=12714 $Y=12936
XX30BB92C5753 GND! VDD! GND! 19 466 228 21 106 227 107 268 
+	269 287 sram_6t $T=12738 12012 0 0 $X=12714 $Y=12012
XX30BB92C5754 GND! VDD! GND! 19 467 229 18 106 225 107 268 
+	269 287 sram_6t $T=14082 12012 0 0 $X=14058 $Y=12012
XX30BB92C5755 GND! VDD! GND! 19 468 230 20 106 226 107 268 
+	269 287 sram_6t $T=13410 12012 0 0 $X=13386 $Y=12012
XX30BB92C5756 GND! VDD! GND! 19 412 231 21 105 228 106 267 
+	268 283 sram_6t $T=12738 11088 0 0 $X=12714 $Y=11088
XX30BB92C5757 GND! VDD! GND! 19 413 232 20 105 230 106 267 
+	268 283 sram_6t $T=13410 11088 0 0 $X=13386 $Y=11088
XX30BB92C5758 GND! VDD! GND! 19 414 233 18 105 229 106 267 
+	268 283 sram_6t $T=14082 11088 0 0 $X=14058 $Y=11088
XX30BB92C5759 GND! VDD! GND! 19 415 234 20 104 232 105 266 
+	267 284 sram_6t $T=13410 10164 0 0 $X=13386 $Y=10164
XX30BB92C5760 GND! VDD! GND! 19 416 235 18 104 233 105 266 
+	267 284 sram_6t $T=14082 10164 0 0 $X=14058 $Y=10164
XX30BB92C5761 GND! VDD! GND! 19 417 236 21 104 231 105 266 
+	267 284 sram_6t $T=12738 10164 0 0 $X=12714 $Y=10164
XX30BB92C5762 GND! VDD! GND! 19 418 164 18 103 235 104 265 
+	266 282 sram_6t $T=14082 9240 0 0 $X=14058 $Y=9240
XX30BB92C5763 GND! VDD! GND! 19 419 162 20 103 234 104 265 
+	266 282 sram_6t $T=13410 9240 0 0 $X=13386 $Y=9240
XX30BB92C5764 GND! VDD! GND! 19 420 160 21 103 236 104 265 
+	266 282 sram_6t $T=12738 9240 0 0 $X=12714 $Y=9240
XX30BB92C5765 GND! VDD! GND! 19 366 159 21 99 160 103 272 
+	265 280 sram_6t $T=12738 8316 0 0 $X=12714 $Y=8316
XX30BB92C5766 GND! VDD! GND! 19 367 161 20 99 162 103 272 
+	265 280 sram_6t $T=13410 8316 0 0 $X=13386 $Y=8316
XX30BB92C5767 GND! VDD! GND! 19 368 163 18 99 164 103 272 
+	265 280 sram_6t $T=14082 8316 0 0 $X=14058 $Y=8316
XX30BB92C5768 GND! VDD! GND! 19 369 501 22 98 157 99 262 
+	272 281 sram_6t $T=14754 7392 0 0 $X=14730 $Y=7392
XX30BB92C5769 GND! VDD! GND! 19 370 502 18 98 163 99 262 
+	272 281 sram_6t $T=14082 7392 0 0 $X=14058 $Y=7392
XX30BB92C5770 GND! VDD! GND! 19 371 495 20 98 161 99 262 
+	272 281 sram_6t $T=13410 7392 0 0 $X=13386 $Y=7392
XX30BB92C5771 GND! VDD! GND! 19 372 496 21 98 159 99 262 
+	272 281 sram_6t $T=12738 7392 0 0 $X=12714 $Y=7392
.ends integration
