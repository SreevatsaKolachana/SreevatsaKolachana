* PEX netlist file	Wed Apr 16 03:43:55 2025	inv
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 0

* Top of hierarchy  cell=inv
.subckt inv GND! VDD! OUT IN 6
*.floating_nets 7 8 9 _GENERATED_10 _GENERATED_11 _GENERATED_12
MM1 OUT IN GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=294  $PIN_XY=252,210,222,294,192,210 $DEVICE_ID=1001
MM2 VDD! IN OUT pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=395  $PIN_XY=420,380,390,395,360,380 $DEVICE_ID=1003
MM3 OUT IN VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=294  $PIN_XY=252,380,222,294,192,380 $DEVICE_ID=1003
.ends inv
