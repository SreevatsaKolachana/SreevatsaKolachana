* PEX netlist file	Thu Apr 17 16:35:22 2025	2to4_decoder_static
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 1
.subckt nor 2 3 4 5 6 7 8 9 10 11 12
.ends nor
.subckt inv 2 3 4 5 6 7 8 10 11 12 13
*.floating_nets 9
.ends inv
.subckt nand 2 3 4 5 6 7 8 11 12 13
*.floating_nets 9 10 14 15
MM1 3 6 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=808 $Y=543  $PIN_XY=838,608,808,543,778,608 $DEVICE_ID=1003
MM2 4 5 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=640 $Y=522  $PIN_XY=670,608,640,522,610,608 $DEVICE_ID=1003
.ends nand
.subckt 2to4_decoder_static_filler_17 2 3 4 5 6 7 8 9
.ends 2to4_decoder_static_filler_17

* Hierarchy Level 0

* Top of hierarchy  cell=2to4_decoder_static
.subckt 2to4_decoder_static VDD! GND! 4 5 6 7 BL0 IN0 OP0 IN0BAR OP0BAR
+	BL1 BL2 BL3 16 17 RS1 19 RS1BAR 21 WS1BAR WS1
+	24 25 26 27 28 29 30 31 WS0BAR RS0BAR 34
+	RS0 WS0 37 38 39 BL0_BAR BL1_BAR BL2_BAR BL3_BAR 52 53
+	54 55 56 57 58 59 60 61 62 63 64
+	65 66 67 68 69 70 71 72 73 74 75
+	76 77 78 79 80 81 82 83
*.floating_nets 89
MM1 IN0BAR 30 BL3_BAR nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2574 $Y=2243  $PIN_XY=2604,2226,2574,2243,2544,2226 $DEVICE_ID=1001
MM2 GND! RS1 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=1197  $PIN_XY=2436,1302,2406,1197,2376,1302 $DEVICE_ID=1001
MM3 39 WS0 116 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=273  $PIN_XY=2436,378,2406,273,2376,378 $DEVICE_ID=1001
MM4 IN0 30 BL3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2238 $Y=2244  $PIN_XY=2268,2226,2238,2244,2208,2226 $DEVICE_ID=1001
MM5 31 17 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2238 $Y=1680  $PIN_XY=2268,1596,2238,1680,2208,1596 $DEVICE_ID=1001
MM6 17 RS0 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=1218  $PIN_XY=2268,1302,2238,1218,2208,1302 $DEVICE_ID=1001
MM7 30 39 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2238 $Y=756  $PIN_XY=2268,672,2238,756,2208,672 $DEVICE_ID=1001
MM8 116 WS1 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=294  $PIN_XY=2268,378,2238,294,2208,378 $DEVICE_ID=1001
MM9 IN0BAR 28 BL2_BAR nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1902 $Y=2243  $PIN_XY=1932,2226,1902,2243,1872,2226 $DEVICE_ID=1001
MM10 GND! RS1 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=1197  $PIN_XY=1764,1302,1734,1197,1704,1302 $DEVICE_ID=1001
MM11 38 WS1 115 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=273  $PIN_XY=1764,378,1734,273,1704,378 $DEVICE_ID=1001
MM12 IN0 28 BL2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1566 $Y=2244  $PIN_XY=1596,2226,1566,2244,1536,2226 $DEVICE_ID=1001
MM13 29 16 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1566 $Y=1680  $PIN_XY=1596,1596,1566,1680,1536,1596 $DEVICE_ID=1001
MM14 16 RS0BAR GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=1218  $PIN_XY=1596,1302,1566,1218,1536,1302 $DEVICE_ID=1001
MM15 28 38 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1566 $Y=756  $PIN_XY=1596,672,1566,756,1536,672 $DEVICE_ID=1001
MM16 115 WS0BAR GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=294  $PIN_XY=1596,378,1566,294,1536,378 $DEVICE_ID=1001
MM17 IN0BAR 26 BL1_BAR nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1230 $Y=2243  $PIN_XY=1260,2226,1230,2243,1200,2226 $DEVICE_ID=1001
MM18 GND! RS1BAR 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=1197  $PIN_XY=1092,1302,1062,1197,1032,1302 $DEVICE_ID=1001
MM19 37 WS0 114 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=273  $PIN_XY=1092,378,1062,273,1032,378 $DEVICE_ID=1001
MM20 IN0 26 BL1 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=894 $Y=2244  $PIN_XY=924,2226,894,2244,864,2226 $DEVICE_ID=1001
MM21 27 19 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=894 $Y=1680  $PIN_XY=924,1596,894,1680,864,1596 $DEVICE_ID=1001
MM22 19 RS0 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=1218  $PIN_XY=924,1302,894,1218,864,1302 $DEVICE_ID=1001
MM23 26 37 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=894 $Y=756  $PIN_XY=924,672,894,756,864,672 $DEVICE_ID=1001
MM24 114 WS1BAR GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=294  $PIN_XY=924,378,894,294,864,378 $DEVICE_ID=1001
MM25 IN0BAR 24 BL0_BAR nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=558 $Y=2243  $PIN_XY=588,2226,558,2243,528,2226 $DEVICE_ID=1001
MM26 GND! RS1BAR 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=1197  $PIN_XY=420,1302,390,1197,360,1302 $DEVICE_ID=1001
MM27 34 WS1BAR 113 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=273  $PIN_XY=420,378,390,273,360,378 $DEVICE_ID=1001
MM28 IN0 24 BL0 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=2267  $PIN_XY=252,2226,222,2267,192,2226 $DEVICE_ID=1001
MM29 25 21 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=1680  $PIN_XY=252,1596,222,1680,192,1596 $DEVICE_ID=1001
MM30 21 RS0BAR GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=1218  $PIN_XY=252,1302,222,1218,192,1302 $DEVICE_ID=1001
MM31 24 34 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=756  $PIN_XY=252,672,222,756,192,672 $DEVICE_ID=1001
MM32 113 WS0BAR GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=294  $PIN_XY=252,378,222,294,192,378 $DEVICE_ID=1001
MM33 OP0BAR 31 BL3_BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2574 $Y=3628  $PIN_XY=2604,3614,2574,3628,2544,3614 $DEVICE_ID=1003
MM34 VDD! 17 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=1781  $PIN_XY=2436,1766,2406,1781,2376,1766 $DEVICE_ID=1003
MM35 17 RS1 112 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=1197  $PIN_XY=2436,1132,2406,1197,2376,1132 $DEVICE_ID=1003
MM36 VDD! 39 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=857  $PIN_XY=2436,842,2406,857,2376,842 $DEVICE_ID=1003
MM37 OP0 31 BL3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2238 $Y=3628  $PIN_XY=2268,3614,2238,3628,2208,3614 $DEVICE_ID=1003
MM38 31 17 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=1680  $PIN_XY=2268,1766,2238,1680,2208,1766 $DEVICE_ID=1003
MM39 112 RS0 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=1218  $PIN_XY=2268,1132,2238,1218,2208,1132 $DEVICE_ID=1003
MM40 30 39 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=756  $PIN_XY=2268,842,2238,756,2208,842 $DEVICE_ID=1003
MM41 OP0BAR 29 BL2_BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1902 $Y=3628  $PIN_XY=1932,3614,1902,3628,1872,3614 $DEVICE_ID=1003
MM42 VDD! 16 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=1781  $PIN_XY=1764,1766,1734,1781,1704,1766 $DEVICE_ID=1003
MM43 16 RS1 111 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=1197  $PIN_XY=1764,1132,1734,1197,1704,1132 $DEVICE_ID=1003
MM44 VDD! 38 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=857  $PIN_XY=1764,842,1734,857,1704,842 $DEVICE_ID=1003
MM45 OP0 29 BL2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1566 $Y=3628  $PIN_XY=1596,3614,1566,3628,1536,3614 $DEVICE_ID=1003
MM46 29 16 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=1680  $PIN_XY=1596,1766,1566,1680,1536,1766 $DEVICE_ID=1003
MM47 111 RS0BAR VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=1218  $PIN_XY=1596,1132,1566,1218,1536,1132 $DEVICE_ID=1003
MM48 28 38 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=756  $PIN_XY=1596,842,1566,756,1536,842 $DEVICE_ID=1003
MM49 OP0BAR 27 BL1_BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1230 $Y=3628  $PIN_XY=1260,3614,1230,3628,1200,3614 $DEVICE_ID=1003
MM50 VDD! 19 27 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=1781  $PIN_XY=1092,1766,1062,1781,1032,1766 $DEVICE_ID=1003
MM51 19 RS1BAR 110 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=1197  $PIN_XY=1092,1132,1062,1197,1032,1132 $DEVICE_ID=1003
MM52 VDD! 37 26 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=857  $PIN_XY=1092,842,1062,857,1032,842 $DEVICE_ID=1003
MM53 OP0 27 BL1 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=894 $Y=3628  $PIN_XY=924,3614,894,3628,864,3614 $DEVICE_ID=1003
MM54 27 19 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=1680  $PIN_XY=924,1766,894,1680,864,1766 $DEVICE_ID=1003
MM55 110 RS0 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=1218  $PIN_XY=924,1132,894,1218,864,1132 $DEVICE_ID=1003
MM56 26 37 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=756  $PIN_XY=924,842,894,756,864,842 $DEVICE_ID=1003
MM57 OP0BAR 25 BL0_BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=558 $Y=3628  $PIN_XY=588,3614,558,3628,528,3614 $DEVICE_ID=1003
MM58 VDD! 21 25 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=1781  $PIN_XY=420,1766,390,1781,360,1766 $DEVICE_ID=1003
MM59 21 RS1BAR 109 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=1197  $PIN_XY=420,1132,390,1197,360,1132 $DEVICE_ID=1003
MM60 VDD! 34 24 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=857  $PIN_XY=420,842,390,857,360,842 $DEVICE_ID=1003
MM61 OP0 25 BL0 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=3628  $PIN_XY=252,3614,222,3628,192,3614 $DEVICE_ID=1003
MM62 25 21 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=1680  $PIN_XY=252,1766,222,1680,192,1766 $DEVICE_ID=1003
MM63 109 RS0BAR VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=1218  $PIN_XY=252,1132,222,1218,192,1132 $DEVICE_ID=1003
MM64 24 34 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=756  $PIN_XY=252,842,222,756,192,842 $DEVICE_ID=1003
XX14806B871 GND! VDD! 29 16 RS0BAR 40 41 84 90 93 101 inv $T=1344 1386 0 0 $X=1344 $Y=1386
XX14806B872 GND! VDD! 31 17 RS0 42 43 84 90 94 102 inv $T=2016 1386 0 0 $X=2016 $Y=1386
XX14806B873 GND! VDD! 27 19 RS0 44 45 84 90 95 103 inv $T=672 1386 0 0 $X=672 $Y=1386
XX14806B874 GND! VDD! 25 21 RS0BAR 46 47 84 90 96 104 inv $T=0 1386 0 0 $X=0 $Y=1386
XX14806B875 GND! VDD! 30 39 WS1 RS0 RS1 85 91 97 105 inv $T=2016 462 0 0 $X=2016 $Y=462
XX14806B876 GND! VDD! 28 38 WS0BAR RS0BAR RS1 85 91 98 106 inv $T=1344 462 0 0 $X=1344 $Y=462
XX14806B877 GND! VDD! 26 37 WS1BAR RS0 RS1BAR 85 91 99 107 inv $T=672 462 0 0 $X=672 $Y=462
XX14806B878 GND! VDD! 24 34 WS0BAR RS0BAR RS1BAR 85 91 100 108 inv $T=0 462 0 0 $X=0 $Y=462
XX14806B879 GND! VDD! _GENERATED_118 VDD! GND! _GENERATED_117 85 92 2to4_decoder_static_filler_17 $T=3132 588 0 180 $X=2688 $Y=-2
XX14806B8710 GND! VDD! GND! _GENERATED_119 _GENERATED_120 VDD! 85 91 2to4_decoder_static_filler_17 $T=2688 462 0 0 $X=2688 $Y=462
XX14806B8711 GND! VDD! _GENERATED_122 VDD! GND! _GENERATED_121 84 91 2to4_decoder_static_filler_17 $T=3132 1512 0 180 $X=2688 $Y=922
XX14806B8712 GND! VDD! GND! _GENERATED_123 _GENERATED_124 VDD! 84 90 2to4_decoder_static_filler_17 $T=2688 1386 0 0 $X=2688 $Y=1386
XX14806B8713 4 VDD! _GENERATED_127 _GENERATED_125 _GENERATED_128 _GENERATED_126 86 90 2to4_decoder_static_filler_17 $T=3132 2436 0 180 $X=2688 $Y=1846
XX14806B8714 4 5 _GENERATED_131 _GENERATED_129 _GENERATED_132 _GENERATED_130 86 BL0 2to4_decoder_static_filler_17 $T=2688 2310 0 0 $X=2688 $Y=2310
XX14806B8715 6 5 _GENERATED_135 _GENERATED_133 _GENERATED_136 _GENERATED_134 87 BL0 2to4_decoder_static_filler_17 $T=3132 3360 0 180 $X=2688 $Y=2770
XX14806B8716 6 7 _GENERATED_139 _GENERATED_137 _GENERATED_140 _GENERATED_138 87 OP0 2to4_decoder_static_filler_17 $T=2688 3234 0 0 $X=2688 $Y=3234
XX14806B8717 GND! VDD! 17 RS1 RS0 17 39 39 112 84 91 nor $T=1388 1514 1 0 $X=2016 $Y=922
XX14806B8718 GND! VDD! 16 RS1 RS0BAR 16 38 38 111 84 91 nor $T=716 1514 1 0 $X=1343 $Y=922
XX14806B8719 GND! VDD! 19 RS1BAR RS0 19 37 37 110 84 91 nor $T=44 1514 1 0 $X=672 $Y=922
XX14806B8720 GND! VDD! 21 RS1BAR RS0BAR 21 34 34 109 84 91 nor $T=-628 1514 1 0 $X=0 $Y=922
XX14806B8721 GND! VDD! 34 WS0BAR WS1BAR 34 113 85 88 92 nand $T=-418 816 1 0 $X=0 $Y=-2
XX14806B8722 GND! VDD! 37 WS1BAR WS0 37 114 85 88 92 nand $T=254 816 1 0 $X=671 $Y=-2
XX14806B8723 GND! VDD! 38 WS0BAR WS1 38 115 85 88 92 nand $T=926 816 1 0 $X=1344 $Y=-2
XX14806B8724 GND! VDD! 39 WS1 WS0 39 116 85 88 92 nand $T=1598 816 1 0 $X=2016 $Y=-2
.ends 2to4_decoder_static
