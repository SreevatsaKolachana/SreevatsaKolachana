* PEX netlist file	Sat Apr 12 17:36:46 2025	nor_layout
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 0

* Top of hierarchy  cell=nor_layout
.subckt nor_layout GND! VDD! Y A B 7 8 9
*.floating_nets 10 11 _GENERATED_12
MM1 GND! B Y nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=478 $Y=522  $PIN_XY=508,438,478,522,448,438 $DEVICE_ID=1001
MM2 Y A GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=142 $Y=522  $PIN_XY=172,438,142,522,112,438 $DEVICE_ID=1001
MM3 VDD! A 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=646 $Y=667  $PIN_XY=676,608,646,667,616,608 $DEVICE_ID=1003
MM4 9 B Y pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=478 $Y=522  $PIN_XY=508,608,478,522,448,608 $DEVICE_ID=1003
MM5 Y B 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=310 $Y=667  $PIN_XY=340,608,310,667,280,608 $DEVICE_ID=1003
MM6 8 A VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=142 $Y=522  $PIN_XY=172,608,142,522,112,608 $DEVICE_ID=1003
.ends nor_layout
