* PEX netlist file	Mon Apr 14 18:18:10 2025	mux_2by1
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 1
.subckt inv 2 3 4 5 7 8 9
*.floating_nets 6 10 11
.ends inv
.subckt nand 2 3 4 5 6 7 8 9 11 12 13
*.floating_nets 10 14 15
MM1 3 6 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=808 $Y=522  $PIN_XY=838,608,808,522,778,608 $DEVICE_ID=1003
MM2 4 5 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=640 $Y=522  $PIN_XY=670,608,640,522,610,608 $DEVICE_ID=1003
.ends nand
.subckt nor 2 3 4 5 6 7 9 10 11
*.floating_nets 12 13 14
MM1 4 6 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1018 $Y=296  $PIN_XY=1048,382,1018,296,988,382 $DEVICE_ID=1003
MM2 8 5 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=850 $Y=296  $PIN_XY=880,382,850,296,820,382 $DEVICE_ID=1003
.ends nor
.subckt sram_filler 2 3 4 5 6
.ends sram_filler

* Hierarchy Level 0

* Top of hierarchy  cell=mux_2by1
.subckt mux_2by1 GND! S 4 5 6 OUT 8
MM1 GND! OUT GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2572 $Y=1384  $PIN_XY=2602,1300,2572,1384,2542,1300 $DEVICE_ID=1001
MM2 GND! 8 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2404 $Y=1384  $PIN_XY=2434,1300,2404,1384,2374,1300 $DEVICE_ID=1001
MM3 16 GND! GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2404 $Y=922  $PIN_XY=2434,1006,2404,922,2374,1006 $DEVICE_ID=1001
MM4 8 6 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1900 $Y=1384  $PIN_XY=1930,1300,1900,1384,1870,1300 $DEVICE_ID=1001
MM5 OUT 5 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1900 $Y=922  $PIN_XY=1930,1006,1900,922,1870,1006 $DEVICE_ID=1001
MM6 6 4 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1396 $Y=1384  $PIN_XY=1426,1300,1396,1384,1366,1300 $DEVICE_ID=1001
MM7 5 10 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1396 $Y=922  $PIN_XY=1426,1006,1396,922,1366,1006 $DEVICE_ID=1001
MM8 18 9 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1228 $Y=1384  $PIN_XY=1258,1300,1228,1384,1198,1300 $DEVICE_ID=1001
MM9 17 S GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1228 $Y=922  $PIN_XY=1258,1006,1228,922,1198,1006 $DEVICE_ID=1001
MM10 4 S GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=724 $Y=1405  $PIN_XY=754,1300,724,1405,694,1300 $DEVICE_ID=1001
MM11 GND! GND! 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2572 $Y=821  $PIN_XY=2602,836,2572,821,2542,836 $DEVICE_ID=1003
MM12 16 GND! GND! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2404 $Y=922  $PIN_XY=2434,836,2404,922,2374,836 $DEVICE_ID=1003
MM13 GND! 6 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2068 $Y=1485  $PIN_XY=2098,1470,2068,1485,2038,1470 $DEVICE_ID=1003
MM14 GND! 5 OUT pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2068 $Y=821  $PIN_XY=2098,836,2068,821,2038,836 $DEVICE_ID=1003
MM15 8 6 GND! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1900 $Y=1384  $PIN_XY=1930,1470,1900,1384,1870,1470 $DEVICE_ID=1003
MM16 OUT 5 GND! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1900 $Y=922  $PIN_XY=1930,836,1900,922,1870,836 $DEVICE_ID=1003
MM17 GND! S 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=892 $Y=1485  $PIN_XY=922,1470,892,1485,862,1470 $DEVICE_ID=1003
MM18 4 S GND! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=724 $Y=1405  $PIN_XY=754,1470,724,1405,694,1470 $DEVICE_ID=1003
XXE8093A5B1 GND! GND! 5 S 10 9 4 17 11 12 14 nand $T=588 1444 1 0 $X=1006 $Y=625
XXE8093A5B2 GND! GND! 6 9 4 S 10 18 11 13 15 nand $T=588 862 0 0 $X=1006 $Y=1090
XXE8093A5B3 GND! GND! 11 13 15 sram_filler $T=2682 1090 0 0 $X=2686 $Y=1090
XXE8093A5B4 GND! GND! 11 12 14 sram_filler $T=3134 1216 0 180 $X=2686 $Y=626
XXE8093A5B5 GND! GND! 11 12 14 sram_filler $T=498 1216 1 0 $X=502 $Y=626
XXE8093A5B6 GND! GND! 11 12 14 sram_filler $T=666 1216 1 0 $X=670 $Y=626
XXE8093A5B7 GND! GND! OUT 5 11 12 14 inv $T=1678 1216 1 0 $X=1678 $Y=626
XXE8093A5B8 GND! GND! 16 GND! 11 12 14 inv $T=2182 1216 1 0 $X=2182 $Y=626
XXE8093A5B9 GND! GND! 8 6 11 13 15 inv $T=1678 1090 0 0 $X=1678 $Y=1090
XXE8093A5B10 GND! GND! 4 S 11 13 15 inv $T=502 1090 0 0 $X=502 $Y=1090
XXE8093A5B11 GND! GND! GND! 8 OUT GND! 11 13 15 nor $T=1554 1088 0 0 $X=2182 $Y=1090
.ends mux_2by1
