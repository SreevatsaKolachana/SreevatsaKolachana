* PEX netlist file	Thu Apr 17 17:21:38 2025	WLRef_PC
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 2
.subckt nor 2 3 4 5 6 7 8 9 10 11
.ends nor
.subckt invx4 2 3 4 5 6 7 8 9 10 11
*.floating_nets 12
.ends invx4
.subckt inv 2 3 4 5 7 8
*.floating_nets 6
.ends inv
.subckt sram_filler 2 3 4 5 6 7
.ends sram_filler
.subckt nand 2 3 4 5 6 7 8 12 13
*.floating_nets 10 11 14 15
MM1 4 6 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=808 $Y=522  $PIN_XY=838,438,808,522,778,438 $DEVICE_ID=1001
MM2 9 5 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=640 $Y=522  $PIN_XY=670,438,640,522,610,438 $DEVICE_ID=1001
.ends nand

* Hierarchy Level 1
.subckt buffer 2 3 4 5 6 7 8
XX5D5DE09B49 2 3 5 4 7 8 inv $T=584 2 0 0 $X=584 $Y=2
XX5D5DE09B50 2 3 4 6 7 8 inv $T=80 2 0 0 $X=80 $Y=2
.ends buffer

* Hierarchy Level 0

* Top of hierarchy  cell=WLRef_PC
.subckt WLRef_PC 9 10 11 12 13 14 15 16 17 18 19
+	20 21 22 23 CLK 25 26 27 28 CLK_DFF 30
+	31 32 33 34 35 WLREF RSNEW PC
*.floating_nets 70 71 72 73 74 75 76 77 78 79 80
*+	81 82 83 84 85 86
MM1 8 35 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5770 $Y=1241  $PIN_XY=5800,1136,5770,1241,5740,1136 $DEVICE_ID=1001
MM2 34 40 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5602 $Y=1661  $PIN_XY=5632,1766,5602,1661,5572,1766 $DEVICE_ID=1001
MM3 35 56 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5602 $Y=737  $PIN_XY=5632,842,5602,737,5572,842 $DEVICE_ID=1001
MM4 8 39 32 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5266 $Y=1241  $PIN_XY=5296,1136,5266,1241,5236,1136 $DEVICE_ID=1001
MM5 40 32 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5098 $Y=1661  $PIN_XY=5128,1766,5098,1661,5068,1766 $DEVICE_ID=1001
MM6 56 30 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5098 $Y=737  $PIN_XY=5128,842,5098,737,5068,842 $DEVICE_ID=1001
MM7 7 27 WLREF nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=2606  $PIN_XY=4792,2690,4762,2606,4732,2690 $DEVICE_ID=1001
MM8 8 31 42 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4762 $Y=1241  $PIN_XY=4792,1136,4762,1241,4732,1136 $DEVICE_ID=1001
MM9 WLREF 27 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4594 $Y=2606  $PIN_XY=4624,2690,4594,2606,4564,2690 $DEVICE_ID=1001
MM10 31 43 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4594 $Y=1682  $PIN_XY=4624,1766,4594,1682,4564,1766 $DEVICE_ID=1001
MM11 30 57 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4594 $Y=737  $PIN_XY=4624,842,4594,737,4564,842 $DEVICE_ID=1001
MM12 4 23 PC nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4426 $Y=2165  $PIN_XY=4456,2060,4426,2165,4396,2060 $DEVICE_ID=1001
MM13 PC 23 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4258 $Y=2165  $PIN_XY=4288,2060,4258,2165,4228,2060 $DEVICE_ID=1001
MM14 8 42 28 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4258 $Y=1241  $PIN_XY=4288,1136,4258,1241,4228,1136 $DEVICE_ID=1001
MM15 43 22 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4090 $Y=1661  $PIN_XY=4120,1766,4090,1661,4060,1766 $DEVICE_ID=1001
MM16 57 28 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4090 $Y=737  $PIN_XY=4120,842,4090,737,4060,842 $DEVICE_ID=1001
MM17 4 12 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3754 $Y=2144  $PIN_XY=3784,2060,3754,2144,3724,2060 $DEVICE_ID=1001
MM18 4 CLK 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3754 $Y=1703  $PIN_XY=3784,1766,3754,1703,3724,1766 $DEVICE_ID=1001
MM19 23 25 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3586 $Y=2165  $PIN_XY=3616,2060,3586,2165,3556,2060 $DEVICE_ID=1001
MM20 4 21 46 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3250 $Y=1661  $PIN_XY=3280,1766,3250,1661,3220,1766 $DEVICE_ID=1001
MM21 8 20 53 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3250 $Y=737  $PIN_XY=3280,842,3250,737,3220,842 $DEVICE_ID=1001
MM22 21 65 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3082 $Y=2144  $PIN_XY=3112,2060,3082,2144,3052,2060 $DEVICE_ID=1001
MM23 20 52 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3082 $Y=1241  $PIN_XY=3112,1136,3082,1241,3052,1136 $DEVICE_ID=1001
MM24 4 46 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2746 $Y=1661  $PIN_XY=2776,1766,2746,1661,2716,1766 $DEVICE_ID=1001
MM25 8 53 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2746 $Y=737  $PIN_XY=2776,842,2746,737,2716,842 $DEVICE_ID=1001
MM26 65 17 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2578 $Y=2144  $PIN_XY=2608,2060,2578,2144,2548,2060 $DEVICE_ID=1001
MM27 52 16 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2578 $Y=1241  $PIN_XY=2608,1136,2578,1241,2548,1136 $DEVICE_ID=1001
MM28 4 19 45 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2242 $Y=1661  $PIN_XY=2272,1766,2242,1661,2212,1766 $DEVICE_ID=1001
MM29 8 18 54 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2242 $Y=737  $PIN_XY=2272,842,2242,737,2212,842 $DEVICE_ID=1001
MM30 17 66 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2074 $Y=2144  $PIN_XY=2104,2060,2074,2144,2044,2060 $DEVICE_ID=1001
MM31 16 51 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2074 $Y=1241  $PIN_XY=2104,1136,2074,1241,2044,1136 $DEVICE_ID=1001
MM32 4 45 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1738 $Y=1661  $PIN_XY=1768,1766,1738,1661,1708,1766 $DEVICE_ID=1001
MM33 8 54 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1738 $Y=737  $PIN_XY=1768,842,1738,737,1708,842 $DEVICE_ID=1001
MM34 66 12 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1570 $Y=2144  $PIN_XY=1600,2060,1570,2144,1540,2060 $DEVICE_ID=1001
MM35 51 11 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1570 $Y=1241  $PIN_XY=1600,1136,1570,1241,1540,1136 $DEVICE_ID=1001
MM36 4 14 44 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1234 $Y=1661  $PIN_XY=1264,1766,1234,1661,1204,1766 $DEVICE_ID=1001
MM37 8 13 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1234 $Y=737  $PIN_XY=1264,842,1234,737,1204,842 $DEVICE_ID=1001
MM38 12 67 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1066 $Y=2144  $PIN_XY=1096,2060,1066,2144,1036,2060 $DEVICE_ID=1001
MM39 11 50 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1066 $Y=1241  $PIN_XY=1096,1136,1066,1241,1036,1136 $DEVICE_ID=1001
MM40 4 44 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=730 $Y=1661  $PIN_XY=760,1766,730,1661,700,1766 $DEVICE_ID=1001
MM41 8 55 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=730 $Y=737  $PIN_XY=760,842,730,737,700,842 $DEVICE_ID=1001
MM42 67 CLK 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=562 $Y=2144  $PIN_XY=592,2060,562,2144,532,2060 $DEVICE_ID=1001
MM43 50 25 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=562 $Y=1241  $PIN_XY=592,1136,562,1241,532,1136 $DEVICE_ID=1001
MM44 3 22 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5602 $Y=296  $PIN_XY=5632,212,5602,296,5572,212 $DEVICE_ID=1001
MM45 33 34 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5434 $Y=275  $PIN_XY=5464,212,5434,275,5404,212 $DEVICE_ID=1001
MM46 3 33 RSNEW nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=296  $PIN_XY=4792,212,4762,296,4732,212 $DEVICE_ID=1001
MM47 RSNEW 33 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4594 $Y=296  $PIN_XY=4624,212,4594,296,4564,212 $DEVICE_ID=1001
MM48 CLK_DFF 41 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4090 $Y=296  $PIN_XY=4120,212,4090,296,4060,212 $DEVICE_ID=1001
MM49 41 26 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3586 $Y=275  $PIN_XY=3616,212,3586,275,3556,212 $DEVICE_ID=1001
MM50 26 49 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3082 $Y=296  $PIN_XY=3112,212,3082,296,3052,212 $DEVICE_ID=1001
MM51 49 15 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2578 $Y=296  $PIN_XY=2608,212,2578,296,2548,212 $DEVICE_ID=1001
MM52 15 48 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2074 $Y=296  $PIN_XY=2104,212,2074,296,2044,212 $DEVICE_ID=1001
MM53 48 10 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1570 $Y=296  $PIN_XY=1600,212,1570,296,1540,212 $DEVICE_ID=1001
MM54 10 47 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1066 $Y=296  $PIN_XY=1096,212,1066,296,1036,212 $DEVICE_ID=1001
MM55 47 9 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=562 $Y=296  $PIN_XY=592,212,562,296,532,212 $DEVICE_ID=1001
MM56 6 40 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5770 $Y=1581  $PIN_XY=5800,1596,5770,1581,5740,1596 $DEVICE_ID=1003
MM57 6 35 39 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5770 $Y=1241  $PIN_XY=5800,1306,5770,1241,5740,1306 $DEVICE_ID=1003
MM58 2 56 35 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5770 $Y=678  $PIN_XY=5800,672,5770,678,5740,672 $DEVICE_ID=1003
MM59 34 40 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5602 $Y=1661  $PIN_XY=5632,1596,5602,1661,5572,1596 $DEVICE_ID=1003
MM60 39 35 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5602 $Y=1321  $PIN_XY=5632,1306,5602,1321,5572,1306 $DEVICE_ID=1003
MM61 35 56 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5602 $Y=737  $PIN_XY=5632,672,5602,737,5572,672 $DEVICE_ID=1003
MM62 6 32 40 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5266 $Y=1581  $PIN_XY=5296,1596,5266,1581,5236,1596 $DEVICE_ID=1003
MM63 6 39 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5266 $Y=1241  $PIN_XY=5296,1306,5266,1241,5236,1306 $DEVICE_ID=1003
MM64 2 30 56 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5266 $Y=678  $PIN_XY=5296,672,5266,678,5236,672 $DEVICE_ID=1003
MM65 40 32 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5098 $Y=1661  $PIN_XY=5128,1596,5098,1661,5068,1596 $DEVICE_ID=1003
MM66 32 39 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5098 $Y=1321  $PIN_XY=5128,1306,5098,1321,5068,1306 $DEVICE_ID=1003
MM67 56 30 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5098 $Y=737  $PIN_XY=5128,672,5098,737,5068,672 $DEVICE_ID=1003
MM68 2 33 RSNEW pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5098 $Y=397  $PIN_XY=5128,382,5098,397,5068,382 $DEVICE_ID=1003
MM69 RSNEW 33 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4930 $Y=376  $PIN_XY=4960,382,4930,376,4900,382 $DEVICE_ID=1003
MM70 5 27 WLREF pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=2606  $PIN_XY=4792,2520,4762,2606,4732,2520 $DEVICE_ID=1003
MM71 5 23 PC pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=2245  $PIN_XY=4792,2230,4762,2245,4732,2230 $DEVICE_ID=1003
MM72 6 43 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=1581  $PIN_XY=4792,1596,4762,1581,4732,1596 $DEVICE_ID=1003
MM73 6 31 42 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=1241  $PIN_XY=4792,1306,4762,1241,4732,1306 $DEVICE_ID=1003
MM74 2 57 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=657  $PIN_XY=4792,672,4762,657,4732,672 $DEVICE_ID=1003
MM75 WLREF 27 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4594 $Y=2606  $PIN_XY=4624,2520,4594,2606,4564,2520 $DEVICE_ID=1003
MM76 PC 23 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4594 $Y=2245  $PIN_XY=4624,2230,4594,2245,4564,2230 $DEVICE_ID=1003
MM77 31 43 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4594 $Y=1682  $PIN_XY=4624,1596,4594,1682,4564,1596 $DEVICE_ID=1003
MM78 42 31 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4594 $Y=1321  $PIN_XY=4624,1306,4594,1321,4564,1306 $DEVICE_ID=1003
MM79 30 57 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4594 $Y=737  $PIN_XY=4624,672,4594,737,4564,672 $DEVICE_ID=1003
MM80 5 27 WLREF pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4426 $Y=2505  $PIN_XY=4456,2520,4426,2505,4396,2520 $DEVICE_ID=1003
MM81 5 23 PC pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4426 $Y=2165  $PIN_XY=4456,2230,4426,2165,4396,2230 $DEVICE_ID=1003
MM82 WLREF 27 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4258 $Y=2505  $PIN_XY=4288,2520,4258,2505,4228,2520 $DEVICE_ID=1003
MM83 PC 23 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4258 $Y=2165  $PIN_XY=4288,2230,4258,2165,4228,2230 $DEVICE_ID=1003
MM84 6 22 43 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4258 $Y=1581  $PIN_XY=4288,1596,4258,1581,4228,1596 $DEVICE_ID=1003
MM85 6 42 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4258 $Y=1241  $PIN_XY=4288,1306,4258,1241,4228,1306 $DEVICE_ID=1003
MM86 2 28 57 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4258 $Y=657  $PIN_XY=4288,672,4258,657,4228,672 $DEVICE_ID=1003
MM87 2 41 CLK_DFF pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4258 $Y=397  $PIN_XY=4288,382,4258,397,4228,382 $DEVICE_ID=1003
MM88 43 22 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4090 $Y=1661  $PIN_XY=4120,1596,4090,1661,4060,1596 $DEVICE_ID=1003
MM89 28 42 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4090 $Y=1321  $PIN_XY=4120,1306,4090,1321,4060,1306 $DEVICE_ID=1003
MM90 57 28 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4090 $Y=737  $PIN_XY=4120,672,4090,737,4060,672 $DEVICE_ID=1003
MM91 5 19 27 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3754 $Y=2606  $PIN_XY=3784,2520,3754,2606,3724,2520 $DEVICE_ID=1003
MM92 23 12 69 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3754 $Y=2144  $PIN_XY=3784,2230,3754,2144,3724,2230 $DEVICE_ID=1003
MM93 6 CLK 22 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3754 $Y=1703  $PIN_XY=3784,1596,3754,1703,3724,1596 $DEVICE_ID=1003
MM94 2 26 41 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3754 $Y=376  $PIN_XY=3784,382,3754,376,3724,382 $DEVICE_ID=1003
MM95 27 12 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3586 $Y=2606  $PIN_XY=3616,2520,3586,2606,3556,2520 $DEVICE_ID=1003
MM96 69 25 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3586 $Y=2165  $PIN_XY=3616,2230,3586,2165,3556,2230 $DEVICE_ID=1003
MM97 22 CLK 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3586 $Y=1602  $PIN_XY=3616,1596,3586,1602,3556,1596 $DEVICE_ID=1003
MM98 5 65 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3250 $Y=2224  $PIN_XY=3280,2230,3250,2224,3220,2230 $DEVICE_ID=1003
MM99 6 21 46 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3250 $Y=1661  $PIN_XY=3280,1596,3250,1661,3220,1596 $DEVICE_ID=1003
MM100 6 52 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3250 $Y=1321  $PIN_XY=3280,1306,3250,1321,3220,1306 $DEVICE_ID=1003
MM101 2 20 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3250 $Y=737  $PIN_XY=3280,672,3250,737,3220,672 $DEVICE_ID=1003
MM102 2 49 26 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3250 $Y=397  $PIN_XY=3280,382,3250,397,3220,382 $DEVICE_ID=1003
MM103 21 65 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3082 $Y=2144  $PIN_XY=3112,2230,3082,2144,3052,2230 $DEVICE_ID=1003
MM104 46 21 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3082 $Y=1581  $PIN_XY=3112,1596,3082,1581,3052,1596 $DEVICE_ID=1003
MM105 20 52 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3082 $Y=1241  $PIN_XY=3112,1306,3082,1241,3052,1306 $DEVICE_ID=1003
MM106 53 20 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3082 $Y=657  $PIN_XY=3112,672,3082,657,3052,672 $DEVICE_ID=1003
MM107 5 17 65 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2746 $Y=2224  $PIN_XY=2776,2230,2746,2224,2716,2230 $DEVICE_ID=1003
MM108 6 46 19 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2746 $Y=1661  $PIN_XY=2776,1596,2746,1661,2716,1596 $DEVICE_ID=1003
MM109 6 16 52 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2746 $Y=1321  $PIN_XY=2776,1306,2746,1321,2716,1306 $DEVICE_ID=1003
MM110 2 53 18 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2746 $Y=737  $PIN_XY=2776,672,2746,737,2716,672 $DEVICE_ID=1003
MM111 2 15 49 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2746 $Y=397  $PIN_XY=2776,382,2746,397,2716,382 $DEVICE_ID=1003
MM112 65 17 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2578 $Y=2144  $PIN_XY=2608,2230,2578,2144,2548,2230 $DEVICE_ID=1003
MM113 19 46 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2578 $Y=1581  $PIN_XY=2608,1596,2578,1581,2548,1596 $DEVICE_ID=1003
MM114 52 16 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2578 $Y=1241  $PIN_XY=2608,1306,2578,1241,2548,1306 $DEVICE_ID=1003
MM115 18 53 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2578 $Y=657  $PIN_XY=2608,672,2578,657,2548,672 $DEVICE_ID=1003
MM116 5 66 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2242 $Y=2224  $PIN_XY=2272,2230,2242,2224,2212,2230 $DEVICE_ID=1003
MM117 6 19 45 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2242 $Y=1661  $PIN_XY=2272,1596,2242,1661,2212,1596 $DEVICE_ID=1003
MM118 6 51 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2242 $Y=1321  $PIN_XY=2272,1306,2242,1321,2212,1306 $DEVICE_ID=1003
MM119 2 18 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2242 $Y=737  $PIN_XY=2272,672,2242,737,2212,672 $DEVICE_ID=1003
MM120 2 48 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2242 $Y=397  $PIN_XY=2272,382,2242,397,2212,382 $DEVICE_ID=1003
MM121 17 66 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2074 $Y=2144  $PIN_XY=2104,2230,2074,2144,2044,2230 $DEVICE_ID=1003
MM122 45 19 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2074 $Y=1581  $PIN_XY=2104,1596,2074,1581,2044,1596 $DEVICE_ID=1003
MM123 16 51 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2074 $Y=1241  $PIN_XY=2104,1306,2074,1241,2044,1306 $DEVICE_ID=1003
MM124 54 18 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2074 $Y=657  $PIN_XY=2104,672,2074,657,2044,672 $DEVICE_ID=1003
MM125 5 12 66 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1738 $Y=2224  $PIN_XY=1768,2230,1738,2224,1708,2230 $DEVICE_ID=1003
MM126 6 45 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1738 $Y=1661  $PIN_XY=1768,1596,1738,1661,1708,1596 $DEVICE_ID=1003
MM127 6 11 51 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1738 $Y=1321  $PIN_XY=1768,1306,1738,1321,1708,1306 $DEVICE_ID=1003
MM128 2 54 13 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1738 $Y=737  $PIN_XY=1768,672,1738,737,1708,672 $DEVICE_ID=1003
MM129 2 10 48 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1738 $Y=397  $PIN_XY=1768,382,1738,397,1708,382 $DEVICE_ID=1003
MM130 66 12 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1570 $Y=2144  $PIN_XY=1600,2230,1570,2144,1540,2230 $DEVICE_ID=1003
MM131 14 45 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1570 $Y=1581  $PIN_XY=1600,1596,1570,1581,1540,1596 $DEVICE_ID=1003
MM132 51 11 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1570 $Y=1241  $PIN_XY=1600,1306,1570,1241,1540,1306 $DEVICE_ID=1003
MM133 13 54 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1570 $Y=657  $PIN_XY=1600,672,1570,657,1540,672 $DEVICE_ID=1003
MM134 5 67 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1234 $Y=2224  $PIN_XY=1264,2230,1234,2224,1204,2230 $DEVICE_ID=1003
MM135 6 14 44 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1234 $Y=1661  $PIN_XY=1264,1596,1234,1661,1204,1596 $DEVICE_ID=1003
MM136 6 50 11 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1234 $Y=1321  $PIN_XY=1264,1306,1234,1321,1204,1306 $DEVICE_ID=1003
MM137 2 13 55 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1234 $Y=737  $PIN_XY=1264,672,1234,737,1204,672 $DEVICE_ID=1003
MM138 2 47 10 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1234 $Y=397  $PIN_XY=1264,382,1234,397,1204,382 $DEVICE_ID=1003
MM139 12 67 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1066 $Y=2144  $PIN_XY=1096,2230,1066,2144,1036,2230 $DEVICE_ID=1003
MM140 44 14 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1066 $Y=1581  $PIN_XY=1096,1596,1066,1581,1036,1596 $DEVICE_ID=1003
MM141 11 50 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1066 $Y=1241  $PIN_XY=1096,1306,1066,1241,1036,1306 $DEVICE_ID=1003
MM142 55 13 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1066 $Y=657  $PIN_XY=1096,672,1066,657,1036,672 $DEVICE_ID=1003
MM143 5 CLK 67 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=730 $Y=2224  $PIN_XY=760,2230,730,2224,700,2230 $DEVICE_ID=1003
MM144 6 44 25 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=730 $Y=1661  $PIN_XY=760,1596,730,1661,700,1596 $DEVICE_ID=1003
MM145 6 25 50 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=730 $Y=1321  $PIN_XY=760,1306,730,1321,700,1306 $DEVICE_ID=1003
MM146 2 55 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=730 $Y=737  $PIN_XY=760,672,730,737,700,672 $DEVICE_ID=1003
MM147 2 9 47 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=730 $Y=397  $PIN_XY=760,382,730,397,700,382 $DEVICE_ID=1003
MM148 67 CLK 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=562 $Y=2144  $PIN_XY=592,2230,562,2144,532,2230 $DEVICE_ID=1003
MM149 25 44 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=562 $Y=1581  $PIN_XY=592,1596,562,1581,532,1596 $DEVICE_ID=1003
MM150 50 25 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=562 $Y=1241  $PIN_XY=592,1306,562,1241,532,1306 $DEVICE_ID=1003
MM151 9 55 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=562 $Y=657  $PIN_XY=592,672,562,657,532,672 $DEVICE_ID=1003
MM152 33 22 68 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5602 $Y=296  $PIN_XY=5632,382,5602,296,5572,382 $DEVICE_ID=1003
MM153 68 34 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5434 $Y=275  $PIN_XY=5464,382,5434,275,5404,382 $DEVICE_ID=1003
MM154 2 33 RSNEW pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4762 $Y=296  $PIN_XY=4792,382,4762,296,4732,382 $DEVICE_ID=1003
MM155 RSNEW 33 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4594 $Y=296  $PIN_XY=4624,382,4594,296,4564,382 $DEVICE_ID=1003
MM156 CLK_DFF 41 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4090 $Y=296  $PIN_XY=4120,382,4090,296,4060,382 $DEVICE_ID=1003
MM157 41 26 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3586 $Y=275  $PIN_XY=3616,382,3586,275,3556,382 $DEVICE_ID=1003
MM158 26 49 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3082 $Y=296  $PIN_XY=3112,382,3082,296,3052,382 $DEVICE_ID=1003
MM159 49 15 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2578 $Y=296  $PIN_XY=2608,382,2578,296,2548,382 $DEVICE_ID=1003
MM160 15 48 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2074 $Y=296  $PIN_XY=2104,382,2074,296,2044,382 $DEVICE_ID=1003
MM161 48 10 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1570 $Y=296  $PIN_XY=1600,382,1570,296,1540,382 $DEVICE_ID=1003
MM162 10 47 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1066 $Y=296  $PIN_XY=1096,382,1066,296,1036,382 $DEVICE_ID=1003
MM163 47 9 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=562 $Y=296  $PIN_XY=592,382,562,296,532,382 $DEVICE_ID=1003
XX5D5DE09B1 3 2 33 22 34 88 56 68 61 62 nor $T=4584 0 0 0 $X=5212 $Y=2
XX5D5DE09B2 4 5 23 12 25 CLK 19 69 59 63 nor $T=2736 1848 0 0 $X=3364 $Y=1850
XX5D5DE09B3 4 6 22 CLK 59 64 inv $T=3976 1976 0 180 $X=3364 $Y=1386
XX5D5DE09B4 7 5 27 12 19 25 12 58 63 nand $T=2946 3128 1 0 $X=3364 $Y=2310
XX5D5DE09B5 8 2 56 35 30 60 62 buffer $T=4796 1054 1 0 $X=4876 $Y=462
XX5D5DE09B6 8 6 39 32 35 60 64 buffer $T=6072 924 1 180 $X=4876 $Y=926
XX5D5DE09B7 4 6 40 34 32 59 64 buffer $T=4796 1978 1 0 $X=4876 $Y=1386
XX5D5DE09B8 3 2 41 CLK_DFF 26 61 62 buffer $T=3284 0 0 0 $X=3364 $Y=2
XX5D5DE09B9 8 2 57 30 28 60 62 buffer $T=3788 1054 1 0 $X=3868 $Y=462
XX5D5DE09B10 8 6 42 28 31 60 64 buffer $T=5064 924 1 180 $X=3868 $Y=926
XX5D5DE09B11 4 6 43 31 22 59 64 buffer $T=3788 1978 1 0 $X=3868 $Y=1386
XX5D5DE09B12 4 6 44 25 14 59 64 buffer $T=1536 1978 0 180 $X=340 $Y=1386
XX5D5DE09B13 4 6 45 14 19 59 64 buffer $T=2544 1978 0 180 $X=1348 $Y=1386
XX5D5DE09B14 4 6 46 19 21 59 64 buffer $T=3552 1978 0 180 $X=2356 $Y=1386
XX5D5DE09B15 4 5 65 21 17 59 63 buffer $T=2276 1848 0 0 $X=2356 $Y=1850
XX5D5DE09B16 4 5 66 17 12 59 63 buffer $T=1268 1848 0 0 $X=1348 $Y=1850
XX5D5DE09B17 4 5 67 12 CLK 59 63 buffer $T=260 1848 0 0 $X=340 $Y=1850
XX5D5DE09B18 3 2 47 10 9 61 62 buffer $T=260 0 0 0 $X=340 $Y=2
XX5D5DE09B19 3 2 48 15 10 61 62 buffer $T=1268 0 0 0 $X=1348 $Y=2
XX5D5DE09B20 3 2 49 26 15 61 62 buffer $T=2276 0 0 0 $X=2356 $Y=2
XX5D5DE09B21 8 6 50 11 25 60 64 buffer $T=260 924 0 0 $X=340 $Y=926
XX5D5DE09B22 8 6 51 16 11 60 64 buffer $T=1268 924 0 0 $X=1348 $Y=926
XX5D5DE09B23 8 6 52 20 16 60 64 buffer $T=2276 924 0 0 $X=2356 $Y=926
XX5D5DE09B24 8 2 53 18 20 60 62 buffer $T=3552 1054 0 180 $X=2356 $Y=462
XX5D5DE09B25 8 2 54 13 18 60 62 buffer $T=2544 1054 0 180 $X=1348 $Y=462
XX5D5DE09B26 8 2 55 9 13 60 62 buffer $T=1536 1054 0 180 $X=340 $Y=462
XX5D5DE09B27 7 5 WLREF 27 23 23 89 23 58 63 invx4 $T=5008 2900 0 180 $X=4035 $Y=2310
XX5D5DE09B28 3 2 RSNEW 33 57 57 87 30 61 62 invx4 $T=4348 2 0 0 $X=4372 $Y=2
XX5D5DE09B29 4 5 PC 23 27 27 43 27 59 63 invx4 $T=4012 1850 0 0 $X=4036 $Y=1850
XX5D5DE09B30 7 5 _GENERATED_91 _GENERATED_90 58 63 sram_filler $T=788 2900 0 180 $X=340 $Y=2310
XX5D5DE09B31 7 5 _GENERATED_93 _GENERATED_92 58 63 sram_filler $T=1124 2900 0 180 $X=676 $Y=2310
XX5D5DE09B32 7 5 _GENERATED_95 _GENERATED_94 58 63 sram_filler $T=1460 2900 0 180 $X=1012 $Y=2310
XX5D5DE09B33 7 5 _GENERATED_97 _GENERATED_96 58 63 sram_filler $T=1796 2900 0 180 $X=1348 $Y=2310
XX5D5DE09B34 7 5 _GENERATED_99 _GENERATED_98 58 63 sram_filler $T=2132 2900 0 180 $X=1684 $Y=2310
XX5D5DE09B35 7 5 _GENERATED_101 _GENERATED_100 58 63 sram_filler $T=2468 2900 0 180 $X=2020 $Y=2310
XX5D5DE09B36 7 5 _GENERATED_103 _GENERATED_102 58 63 sram_filler $T=2804 2900 0 180 $X=2356 $Y=2310
XX5D5DE09B37 7 5 _GENERATED_105 _GENERATED_104 58 63 sram_filler $T=3140 2900 0 180 $X=2692 $Y=2310
XX5D5DE09B38 7 5 _GENERATED_107 _GENERATED_106 58 63 sram_filler $T=3476 2900 0 180 $X=3028 $Y=2310
XX5D5DE09B39 7 5 _GENERATED_109 _GENERATED_108 58 63 sram_filler $T=5996 2900 0 180 $X=5548 $Y=2310
XX5D5DE09B40 7 5 _GENERATED_111 _GENERATED_110 58 63 sram_filler $T=5660 2900 0 180 $X=5212 $Y=2310
XX5D5DE09B41 7 5 _GENERATED_113 _GENERATED_112 58 63 sram_filler $T=5324 2900 0 180 $X=4875 $Y=2310
XX5D5DE09B42 4 5 _GENERATED_115 _GENERATED_114 59 63 sram_filler $T=5544 1850 0 0 $X=5548 $Y=1850
XX5D5DE09B43 4 5 _GENERATED_117 _GENERATED_116 59 63 sram_filler $T=5208 1850 0 0 $X=5212 $Y=1850
XX5D5DE09B44 4 5 _GENERATED_119 _GENERATED_118 59 63 sram_filler $T=4872 1850 0 0 $X=4875 $Y=1850
XX5D5DE09B45 8 2 2 _GENERATED_120 60 62 sram_filler $T=3812 1052 0 180 $X=3364 $Y=462
XX5D5DE09B46 8 2 _GENERATED_121 8 60 62 sram_filler $T=3980 1052 0 180 $X=3532 $Y=462
XX5D5DE09B47 8 6 6 _GENERATED_122 60 64 sram_filler $T=3528 926 0 0 $X=3532 $Y=926
XX5D5DE09B48 8 6 _GENERATED_123 8 60 64 sram_filler $T=3360 926 0 0 $X=3364 $Y=926
.ends WLRef_PC
