* PEX netlist file	Tue Apr 15 19:38:09 2025	Demux
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 1
.subckt inv 2 3 4 5 7 8 9
*.floating_nets 6 10 11
.ends inv
.subckt nand 2 3 4 5 6 7 8 9 12 13 14
*.floating_nets 10 11 15 16
MM1 3 6 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=808 $Y=522  $PIN_XY=838,608,808,522,778,608 $DEVICE_ID=1003
MM2 4 5 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=640 $Y=522  $PIN_XY=670,608,640,522,610,608 $DEVICE_ID=1003
.ends nand
.subckt sram_filler 2 3 4 5 6 7 8
.ends sram_filler

* Hierarchy Level 0

* Top of hierarchy  cell=Demux
.subckt Demux VDD! GND! SEL 5 A Y1 Y0
MM1 15 Y0 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1398 $Y=756  $PIN_XY=1428,672,1398,756,1368,672 $DEVICE_ID=1001
MM2 14 Y1 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1398 $Y=294  $PIN_XY=1428,378,1398,294,1368,378 $DEVICE_ID=1001
MM3 Y0 5 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=894 $Y=756  $PIN_XY=924,672,894,756,864,672 $DEVICE_ID=1001
MM4 Y1 SEL 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=894 $Y=294  $PIN_XY=924,378,894,294,864,378 $DEVICE_ID=1001
MM5 17 A GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=726 $Y=756  $PIN_XY=756,672,726,756,696,672 $DEVICE_ID=1001
MM6 16 A GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=726 $Y=294  $PIN_XY=756,378,726,294,696,378 $DEVICE_ID=1001
MM7 5 SEL GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=777  $PIN_XY=252,672,222,777,192,672 $DEVICE_ID=1001
MM8 VDD! Y0 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1566 $Y=857  $PIN_XY=1596,842,1566,857,1536,842 $DEVICE_ID=1003
MM9 VDD! Y1 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1566 $Y=193  $PIN_XY=1596,208,1566,193,1536,208 $DEVICE_ID=1003
MM10 15 Y0 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1398 $Y=756  $PIN_XY=1428,842,1398,756,1368,842 $DEVICE_ID=1003
MM11 14 Y1 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1398 $Y=294  $PIN_XY=1428,208,1398,294,1368,208 $DEVICE_ID=1003
MM12 VDD! SEL 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=857  $PIN_XY=420,842,390,857,360,842 $DEVICE_ID=1003
MM13 5 SEL VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=777  $PIN_XY=252,842,222,777,192,842 $DEVICE_ID=1003
XXACF9D7931 GND! VDD! Y0 A 5 A SEL 17 9 10 12 nand $T=86 234 0 0 $X=504 $Y=462
XXACF9D7932 GND! VDD! Y1 A SEL A 5 16 9 11 13 nand $T=86 816 1 0 $X=504 $Y=-2
XXACF9D7933 GND! VDD! 5 SEL 9 10 12 inv $T=0 462 0 0 $X=0 $Y=462
XXACF9D7934 GND! VDD! 15 Y0 9 10 12 inv $T=1176 462 0 0 $X=1176 $Y=462
XXACF9D7935 GND! VDD! 14 Y1 9 11 13 inv $T=1176 588 1 0 $X=1176 $Y=-2
XXACF9D7936 GND! VDD! _GENERATED_18 GND! 9 11 13 sram_filler $T=616 588 0 180 $X=167 $Y=-2
XXACF9D7937 GND! VDD! VDD! _GENERATED_19 9 11 13 sram_filler $T=448 588 0 180 $X=0 $Y=-2
XXACF9D7938 GND! VDD! _GENERATED_21 _GENERATED_20 9 10 12 sram_filler $T=1676 462 0 0 $X=1680 $Y=462
XXACF9D7939 GND! VDD! VDD! _GENERATED_22 9 11 13 sram_filler $T=2128 588 0 180 $X=1680 $Y=-2
.ends Demux
