* PEX netlist file	Tue Apr 15 19:47:28 2025	buffer_highdrive_vertical
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 1
.subckt invx4 2 3 4 5 6 7 8 9 10
*.floating_nets 11 12 13 14
MM1 3 5 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=750 $Y=395  $PIN_XY=780,380,750,395,720,380 $DEVICE_ID=1003
MM2 4 5 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=582 $Y=395  $PIN_XY=612,380,582,395,552,380 $DEVICE_ID=1003
MM3 3 5 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=414 $Y=294  $PIN_XY=444,380,414,294,384,380 $DEVICE_ID=1003
MM4 4 5 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=246 $Y=294  $PIN_XY=276,380,246,294,216,380 $DEVICE_ID=1003
.ends invx4
.subckt sram_filler 2 3 6 7 8
*.floating_nets 4 5
.ends sram_filler

* Hierarchy Level 0

* Top of hierarchy  cell=buffer_highdrive_vertical
.subckt buffer_highdrive_vertical GND! VDD! 4 OUT IN
MM1 GND! IN 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=392 $Y=292  $PIN_XY=422,208,392,292,362,208 $DEVICE_ID=1001
MM2 GND! 4 OUT nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=392 $Y=-170  $PIN_XY=422,-86,392,-170,362,-86 $DEVICE_ID=1001
MM3 4 IN GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=224 $Y=292  $PIN_XY=254,208,224,292,194,208 $DEVICE_ID=1001
MM4 OUT 4 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=224 $Y=-170  $PIN_XY=254,-86,224,-170,194,-86 $DEVICE_ID=1001
XXBDB3BE301 GND! VDD! 7 8 10 sram_filler $T=838 -2 0 0 $X=842 $Y=-2
XXBDB3BE302 GND! VDD! 7 9 11 sram_filler $T=838 124 1 0 $X=842 $Y=-465
XXBDB3BE303 GND! VDD! 4 IN 4 4 7 8 10 invx4 $T=-22 -2 0 0 $X=2 $Y=-2
XXBDB3BE304 GND! VDD! OUT 4 IN IN 7 9 11 invx4 $T=-22 124 1 0 $X=2 $Y=-465
.ends buffer_highdrive_vertical
