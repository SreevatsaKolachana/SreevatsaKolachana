* PEX netlist file	Thu Apr 17 00:00:55 2025	between_blocks
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 1
.subckt nor 2 3 4 5 6 7 8 9 10 11
.ends nor
.subckt inv 2 3 4 5 6 7 9 10
*.floating_nets 8
.ends inv
.subckt nand 2 3 4 5 6 7 8 9 12 13
*.floating_nets 10 11
.ends nand
.subckt sram_filler 2 3 6 7
*.floating_nets 4 5
.ends sram_filler

* Hierarchy Level 0

* Top of hierarchy  cell=between_blocks
.subckt between_blocks GND! VDD! 4 5 6 7 RSNEW WLREF RS1BAR RS1 RS0
+	RS0BAR 14 15 16 17
*.floating_nets 43 44 _GENERATED_287 _GENERATED_288
MM1 GND! 15 41 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1390 $Y=1777  $PIN_XY=1420,1882,1390,1777,1360,1882 $DEVICE_ID=1001
MM2 GND! 14 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1390 $Y=853  $PIN_XY=1420,958,1390,853,1360,958 $DEVICE_ID=1001
MM3 GND! 7 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1390 $Y=-71  $PIN_XY=1420,34,1390,-71,1360,34 $DEVICE_ID=1001
MM4 GND! 6 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1390 $Y=-995  $PIN_XY=1420,-890,1390,-995,1360,-890 $DEVICE_ID=1001
MM5 42 5 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1222 $Y=2281  $PIN_XY=1252,2176,1222,2281,1192,2176 $DEVICE_ID=1001
MM6 40 4 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1222 $Y=1357  $PIN_XY=1252,1252,1222,1357,1192,1252 $DEVICE_ID=1001
MM7 38 17 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1222 $Y=433  $PIN_XY=1252,328,1222,433,1192,328 $DEVICE_ID=1001
MM8 36 16 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1222 $Y=-491  $PIN_XY=1252,-596,1222,-491,1192,-596 $DEVICE_ID=1001
MM9 GND! RSNEW 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=1798  $PIN_XY=916,1882,886,1798,856,1882 $DEVICE_ID=1001
MM10 GND! RSNEW 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=874  $PIN_XY=916,958,886,874,856,958 $DEVICE_ID=1001
MM11 GND! WLREF 34 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=-50  $PIN_XY=916,34,886,-50,856,34 $DEVICE_ID=1001
MM12 GND! WLREF 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=-995  $PIN_XY=916,-890,886,-995,856,-890 $DEVICE_ID=1001
MM13 GND! RS0 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=2260  $PIN_XY=748,2176,718,2260,688,2176 $DEVICE_ID=1001
MM14 15 RS0BAR GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=1798  $PIN_XY=748,1882,718,1798,688,1882 $DEVICE_ID=1001
MM15 GND! RS1 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=1336  $PIN_XY=748,1252,718,1336,688,1252 $DEVICE_ID=1001
MM16 14 RS1BAR GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=874  $PIN_XY=748,958,718,874,688,958 $DEVICE_ID=1001
MM17 17 18 32 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=412  $PIN_XY=748,328,718,412,688,328 $DEVICE_ID=1001
MM18 34 21 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=-50  $PIN_XY=748,34,718,-50,688,34 $DEVICE_ID=1001
MM19 16 19 31 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=-512  $PIN_XY=748,-596,718,-512,688,-596 $DEVICE_ID=1001
MM20 33 20 6 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=-974  $PIN_XY=748,-890,718,-974,688,-890 $DEVICE_ID=1001
MM21 5 RSNEW GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=2281  $PIN_XY=580,2176,550,2281,520,2176 $DEVICE_ID=1001
MM22 4 RSNEW GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=1336  $PIN_XY=580,1252,550,1336,520,1252 $DEVICE_ID=1001
MM23 32 WLREF GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=412  $PIN_XY=580,328,550,412,520,328 $DEVICE_ID=1001
MM24 31 WLREF GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=-512  $PIN_XY=580,-596,550,-512,520,-596 $DEVICE_ID=1001
MM25 VDD! 5 42 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=2361  $PIN_XY=1420,2346,1390,2361,1360,2346 $DEVICE_ID=1003
MM26 VDD! 15 41 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=1777  $PIN_XY=1420,1712,1390,1777,1360,1712 $DEVICE_ID=1003
MM27 VDD! 4 40 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=1437  $PIN_XY=1420,1422,1390,1437,1360,1422 $DEVICE_ID=1003
MM28 VDD! 14 39 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=853  $PIN_XY=1420,788,1390,853,1360,788 $DEVICE_ID=1003
MM29 VDD! 17 38 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=513  $PIN_XY=1420,498,1390,513,1360,498 $DEVICE_ID=1003
MM30 VDD! 7 37 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=-71  $PIN_XY=1420,-136,1390,-71,1360,-136 $DEVICE_ID=1003
MM31 VDD! 16 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=-411  $PIN_XY=1420,-426,1390,-411,1360,-426 $DEVICE_ID=1003
MM32 VDD! 6 35 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=-995  $PIN_XY=1420,-1060,1390,-995,1360,-1060 $DEVICE_ID=1003
MM33 42 5 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=2281  $PIN_XY=1252,2346,1222,2281,1192,2346 $DEVICE_ID=1003
MM34 41 15 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=1697  $PIN_XY=1252,1712,1222,1697,1192,1712 $DEVICE_ID=1003
MM35 40 4 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=1357  $PIN_XY=1252,1422,1222,1357,1192,1422 $DEVICE_ID=1003
MM36 39 14 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=773  $PIN_XY=1252,788,1222,773,1192,788 $DEVICE_ID=1003
MM37 38 17 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=433  $PIN_XY=1252,498,1222,433,1192,498 $DEVICE_ID=1003
MM38 37 7 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=-151  $PIN_XY=1252,-136,1222,-151,1192,-136 $DEVICE_ID=1003
MM39 36 16 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=-491  $PIN_XY=1252,-426,1222,-491,1192,-426 $DEVICE_ID=1003
MM40 35 6 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=-1075  $PIN_XY=1252,-1060,1222,-1075,1192,-1060 $DEVICE_ID=1003
MM41 VDD! RSNEW 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=1798  $PIN_XY=916,1712,886,1798,856,1712 $DEVICE_ID=1003
MM42 VDD! RSNEW 51 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=874  $PIN_XY=916,788,886,874,856,788 $DEVICE_ID=1003
MM43 VDD! WLREF 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=-50  $PIN_XY=916,-136,886,-50,856,-136 $DEVICE_ID=1003
MM44 VDD! WLREF 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=-995  $PIN_XY=916,-1060,886,-995,856,-1060 $DEVICE_ID=1003
MM45 5 RS0 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=2260  $PIN_XY=748,2346,718,2260,688,2346 $DEVICE_ID=1003
MM46 53 RS0BAR 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=1798  $PIN_XY=748,1712,718,1798,688,1712 $DEVICE_ID=1003
MM47 4 RS1 52 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=1336  $PIN_XY=748,1422,718,1336,688,1422 $DEVICE_ID=1003
MM48 51 RS1BAR 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=874  $PIN_XY=748,788,718,874,688,788 $DEVICE_ID=1003
MM49 VDD! 18 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=412  $PIN_XY=748,498,718,412,688,498 $DEVICE_ID=1003
MM50 7 21 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=-50  $PIN_XY=748,-136,718,-50,688,-136 $DEVICE_ID=1003
MM51 VDD! 19 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=-512  $PIN_XY=748,-426,718,-512,688,-426 $DEVICE_ID=1003
MM52 6 20 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=-974  $PIN_XY=748,-1060,718,-974,688,-1060 $DEVICE_ID=1003
MM53 54 RSNEW VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=2281  $PIN_XY=580,2346,550,2281,520,2346 $DEVICE_ID=1003
MM54 52 RSNEW VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=1336  $PIN_XY=580,1422,550,1336,520,1422 $DEVICE_ID=1003
MM55 17 WLREF VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=412  $PIN_XY=580,498,550,412,520,498 $DEVICE_ID=1003
MM56 16 WLREF VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=-512  $PIN_XY=580,-426,550,-512,520,-426 $DEVICE_ID=1003
XX30C0E9261 GND! VDD! 35 6 49 47 22 26 inv $T=1612 -680 0 180 $X=1000 $Y=-1270
XX30C0E9262 GND! VDD! 36 16 7 7 22 27 inv $T=1000 -806 0 0 $X=1000 $Y=-806
XX30C0E9263 GND! VDD! 37 7 16 16 23 27 inv $T=1612 244 0 180 $X=1000 $Y=-346
XX30C0E9264 GND! VDD! 38 17 14 14 23 28 inv $T=1000 118 0 0 $X=1000 $Y=118
XX30C0E9265 GND! VDD! 39 14 17 17 24 28 inv $T=1612 1168 0 180 $X=1000 $Y=578
XX30C0E9266 GND! VDD! 40 4 15 15 24 29 inv $T=1000 1042 0 0 $X=1000 $Y=1042
XX30C0E9267 GND! VDD! 41 15 4 4 25 29 inv $T=1612 2092 0 180 $X=1000 $Y=1502
XX30C0E9268 GND! VDD! 42 5 48 50 25 30 inv $T=1000 1966 0 0 $X=1000 $Y=1966
XX30C0E9269 GND! VDD! 22 26 sram_filler $T=1952 -680 0 180 $X=1504 $Y=-1270
XX30C0E92610 GND! VDD! 22 27 sram_filler $T=1500 -806 0 0 $X=1504 $Y=-806
XX30C0E92611 GND! VDD! 23 27 sram_filler $T=1952 244 0 180 $X=1504 $Y=-346
XX30C0E92612 GND! VDD! 23 28 sram_filler $T=1500 118 0 0 $X=1504 $Y=118
XX30C0E92613 GND! VDD! 24 28 sram_filler $T=1952 1168 0 180 $X=1504 $Y=578
XX30C0E92614 GND! VDD! 24 29 sram_filler $T=1500 1042 0 0 $X=1504 $Y=1042
XX30C0E92615 GND! VDD! 25 29 sram_filler $T=1952 2092 0 180 $X=1504 $Y=1502
XX30C0E92616 GND! VDD! 25 30 sram_filler $T=1500 1966 0 0 $X=1504 $Y=1966
XX30C0E92617 GND! VDD! 14 RSNEW RS1BAR RS1 18 51 24 28 nor $T=1736 1170 0 180 $X=328 $Y=578
XX30C0E92618 GND! VDD! 4 RSNEW RS1 RS1BAR RS0BAR 52 24 29 nor $T=-300 1040 0 0 $X=328 $Y=1042
XX30C0E92619 GND! VDD! 15 RSNEW RS0BAR RS0 RS1 53 25 29 nor $T=1736 2094 0 180 $X=328 $Y=1501
XX30C0E92620 GND! VDD! 5 RSNEW RS0 RS0BAR 46 54 25 30 nor $T=-300 1964 0 0 $X=328 $Y=1966
XX30C0E92621 GND! VDD! 6 WLREF 20 19 45 33 22 26 nand $T=1526 -452 0 180 $X=328 $Y=-1270
XX30C0E92622 GND! VDD! 16 WLREF 19 20 21 31 22 27 nand $T=-90 -1034 0 0 $X=327 $Y=-806
XX30C0E92623 GND! VDD! 7 WLREF 21 18 19 34 23 27 nand $T=1526 472 0 180 $X=328 $Y=-346
XX30C0E92624 GND! VDD! 17 WLREF 18 21 RS1BAR 32 23 28 nand $T=-90 -110 0 0 $X=327 $Y=118
.ends between_blocks
