* PEX netlist file	Fri Apr 18 05:52:32 2025	memory_array_static_column_decoder_test
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 3
.subckt sram_filler 2 3 4 5 6 7
.ends sram_filler
.subckt tspc_pos_ff 2 3 4 8 9 25 26 27
*.floating_nets 10 11 13 14 15 17 18 19 20 22 23
*+	24 28 29 30 31 32 33 34 35
MM1 4 7 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1176 $Y=294  $PIN_XY=1206,210,1176,294,1146,210 $DEVICE_ID=1001
MM2 2 6 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1008 $Y=294  $PIN_XY=1038,210,1008,294,978,210 $DEVICE_ID=1001
MM3 16 9 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=840 $Y=209  $PIN_XY=870,210,840,209,810,210 $DEVICE_ID=1001
MM4 6 9 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=504 $Y=209  $PIN_XY=534,210,504,209,474,210 $DEVICE_ID=1001
MM5 12 5 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=336 $Y=209  $PIN_XY=366,210,336,209,306,210 $DEVICE_ID=1001
MM6 2 8 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=168 $Y=209  $PIN_XY=198,210,168,209,138,210 $DEVICE_ID=1001
MM7 4 7 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1176 $Y=294  $PIN_XY=1206,380,1176,294,1146,380 $DEVICE_ID=1003
MM8 3 6 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1008 $Y=294  $PIN_XY=1038,380,1008,294,978,380 $DEVICE_ID=1003
MM9 5 9 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=504 $Y=649  $PIN_XY=534,670,504,649,474,670 $DEVICE_ID=1003
MM10 21 8 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=336 $Y=670  $PIN_XY=366,670,336,670,306,670 $DEVICE_ID=1003
MM11 3 9 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=168 $Y=670  $PIN_XY=198,670,168,670,138,670 $DEVICE_ID=1003
.ends tspc_pos_ff
.subckt nand 2 3 4 5 6 7 10 11
*.floating_nets 8 9
.ends nand
.subckt inv 2 3 4 5 7 8
*.floating_nets 6
.ends inv
.subckt 2to4_decoder_static_filler_17 2 3 4 5 6 7
.ends 2to4_decoder_static_filler_17
.subckt Filler 2 3 4 5 6 7 8 9
.ends Filler
.subckt precharge_logic 2 3 4 5 6 7 8 11 12
*.floating_nets 9 10
.ends precharge_logic
.subckt sram_6t 2 3 4 5 6 7 8 9 10 11 14
+	15 16
*.floating_nets 12 13 17 18
MM1 3 6 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=366 $Y=756  $PIN_XY=396,670,366,756,336,670 $DEVICE_ID=1003
.ends sram_6t
.subckt bitcell_precharge_filler 2 3 4 5 6 7
.ends bitcell_precharge_filler
.subckt nor 2 3 4 5 6 7 8 9
.ends nor
.subckt invx4 2 3 4 5 6 7
.ends invx4

* Hierarchy Level 2
.subckt 2to4_decoder_static 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16 17 18 19 20 21 22 25
+	27 29 30 32 34 36 38 39 40 41 42
+	43 44 45 46 79 80 81 82 83 84 85
+	86 87
*.floating_nets 47 48 49 50 51 52 53 54 55 56 57
*+	58 59 60 61 62 63 64 65 66 67 68
*+	69 70 71 72 73 74 75 76 77 78 96
*+	97 98 99 100 101 102 103
MM1 21 37 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2574 $Y=2243  $PIN_XY=2604,2226,2574,2243,2544,2226 $DEVICE_ID=1001
MM2 5 25 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=1197  $PIN_XY=2436,1302,2406,1197,2376,1302 $DEVICE_ID=1001
MM3 46 43 95 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=294  $PIN_XY=2436,378,2406,294,2376,378 $DEVICE_ID=1001
MM4 17 37 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2238 $Y=2244  $PIN_XY=2268,2226,2238,2244,2208,2226 $DEVICE_ID=1001
MM5 38 24 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2238 $Y=1680  $PIN_XY=2268,1596,2238,1680,2208,1596 $DEVICE_ID=1001
MM6 24 42 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=1218  $PIN_XY=2268,1302,2238,1218,2208,1302 $DEVICE_ID=1001
MM7 37 46 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2238 $Y=756  $PIN_XY=2268,672,2238,756,2208,672 $DEVICE_ID=1001
MM8 95 30 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=315  $PIN_XY=2268,378,2238,315,2208,378 $DEVICE_ID=1001
MM9 21 35 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1902 $Y=2243  $PIN_XY=1932,2226,1902,2243,1872,2226 $DEVICE_ID=1001
MM10 5 25 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=1197  $PIN_XY=1764,1302,1734,1197,1704,1302 $DEVICE_ID=1001
MM11 45 30 94 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=294  $PIN_XY=1764,378,1734,294,1704,378 $DEVICE_ID=1001
MM12 15 35 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1566 $Y=2244  $PIN_XY=1596,2226,1566,2244,1536,2226 $DEVICE_ID=1001
MM13 36 23 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1566 $Y=1680  $PIN_XY=1596,1596,1566,1680,1536,1596 $DEVICE_ID=1001
MM14 23 40 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=1218  $PIN_XY=1596,1302,1566,1218,1536,1302 $DEVICE_ID=1001
MM15 35 45 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1566 $Y=756  $PIN_XY=1596,672,1566,756,1536,672 $DEVICE_ID=1001
MM16 94 39 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=315  $PIN_XY=1596,378,1566,315,1536,378 $DEVICE_ID=1001
MM17 21 33 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1230 $Y=2243  $PIN_XY=1260,2226,1230,2243,1200,2226 $DEVICE_ID=1001
MM18 5 27 26 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=1197  $PIN_XY=1092,1302,1062,1197,1032,1302 $DEVICE_ID=1001
MM19 44 43 93 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=294  $PIN_XY=1092,378,1062,294,1032,378 $DEVICE_ID=1001
MM20 13 33 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=894 $Y=2244  $PIN_XY=924,2226,894,2244,864,2226 $DEVICE_ID=1001
MM21 34 26 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=894 $Y=1680  $PIN_XY=924,1596,894,1680,864,1596 $DEVICE_ID=1001
MM22 26 42 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=1218  $PIN_XY=924,1302,894,1218,864,1302 $DEVICE_ID=1001
MM23 33 44 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=894 $Y=756  $PIN_XY=924,672,894,756,864,672 $DEVICE_ID=1001
MM24 93 29 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=315  $PIN_XY=924,378,894,315,864,378 $DEVICE_ID=1001
MM25 21 31 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=558 $Y=2243  $PIN_XY=588,2226,558,2243,528,2226 $DEVICE_ID=1001
MM26 5 27 28 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=1197  $PIN_XY=420,1302,390,1197,360,1302 $DEVICE_ID=1001
MM27 41 29 92 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=294  $PIN_XY=420,378,390,294,360,378 $DEVICE_ID=1001
MM28 11 31 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=2267  $PIN_XY=252,2226,222,2267,192,2226 $DEVICE_ID=1001
MM29 32 28 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=1680  $PIN_XY=252,1596,222,1680,192,1596 $DEVICE_ID=1001
MM30 28 40 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=1218  $PIN_XY=252,1302,222,1218,192,1302 $DEVICE_ID=1001
MM31 31 41 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=756  $PIN_XY=252,672,222,756,192,672 $DEVICE_ID=1001
MM32 92 39 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=315  $PIN_XY=252,378,222,315,192,378 $DEVICE_ID=1001
MM33 6 24 38 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=1781  $PIN_XY=2436,1766,2406,1781,2376,1766 $DEVICE_ID=1003
MM34 24 25 88 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=1197  $PIN_XY=2436,1132,2406,1197,2376,1132 $DEVICE_ID=1003
MM35 4 46 37 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=857  $PIN_XY=2436,842,2406,857,2376,842 $DEVICE_ID=1003
MM36 38 24 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=1680  $PIN_XY=2268,1766,2238,1680,2208,1766 $DEVICE_ID=1003
MM37 88 42 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=1218  $PIN_XY=2268,1132,2238,1218,2208,1132 $DEVICE_ID=1003
MM38 37 46 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=756  $PIN_XY=2268,842,2238,756,2208,842 $DEVICE_ID=1003
MM39 6 23 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=1781  $PIN_XY=1764,1766,1734,1781,1704,1766 $DEVICE_ID=1003
MM40 23 25 89 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=1197  $PIN_XY=1764,1132,1734,1197,1704,1132 $DEVICE_ID=1003
MM41 4 45 35 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=857  $PIN_XY=1764,842,1734,857,1704,842 $DEVICE_ID=1003
MM42 36 23 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=1680  $PIN_XY=1596,1766,1566,1680,1536,1766 $DEVICE_ID=1003
MM43 89 40 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=1218  $PIN_XY=1596,1132,1566,1218,1536,1132 $DEVICE_ID=1003
MM44 35 45 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=756  $PIN_XY=1596,842,1566,756,1536,842 $DEVICE_ID=1003
MM45 6 26 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=1781  $PIN_XY=1092,1766,1062,1781,1032,1766 $DEVICE_ID=1003
MM46 26 27 90 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=1197  $PIN_XY=1092,1132,1062,1197,1032,1132 $DEVICE_ID=1003
MM47 4 44 33 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=857  $PIN_XY=1092,842,1062,857,1032,842 $DEVICE_ID=1003
MM48 34 26 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=1680  $PIN_XY=924,1766,894,1680,864,1766 $DEVICE_ID=1003
MM49 90 42 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=1218  $PIN_XY=924,1132,894,1218,864,1132 $DEVICE_ID=1003
MM50 33 44 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=756  $PIN_XY=924,842,894,756,864,842 $DEVICE_ID=1003
MM51 6 28 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=1781  $PIN_XY=420,1766,390,1781,360,1766 $DEVICE_ID=1003
MM52 28 27 91 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=1197  $PIN_XY=420,1132,390,1197,360,1132 $DEVICE_ID=1003
MM53 4 41 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=857  $PIN_XY=420,842,390,857,360,842 $DEVICE_ID=1003
MM54 32 28 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=1680  $PIN_XY=252,1766,222,1680,192,1766 $DEVICE_ID=1003
MM55 91 40 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=1218  $PIN_XY=252,1132,222,1218,192,1132 $DEVICE_ID=1003
MM56 31 41 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=756  $PIN_XY=252,842,222,756,192,842 $DEVICE_ID=1003
XXB19A871F999 5 6 36 23 79 83 inv $T=1344 1386 0 0 $X=1344 $Y=1386
XXB19A871F1000 5 6 38 24 79 83 inv $T=2016 1386 0 0 $X=2016 $Y=1386
XXB19A871F1001 5 6 34 26 79 83 inv $T=672 1386 0 0 $X=672 $Y=1386
XXB19A871F1002 5 6 32 28 79 83 inv $T=0 1386 0 0 $X=0 $Y=1386
XXB19A871F1003 3 4 37 46 80 84 inv $T=2016 462 0 0 $X=2016 $Y=462
XXB19A871F1004 3 4 35 45 80 84 inv $T=1344 462 0 0 $X=1344 $Y=462
XXB19A871F1005 3 4 33 44 80 84 inv $T=672 462 0 0 $X=672 $Y=462
XXB19A871F1006 3 4 31 41 80 84 inv $T=0 462 0 0 $X=0 $Y=462
XXB19A871F1007 5 4 24 25 42 88 79 84 nor $T=1388 1514 1 0 $X=2016 $Y=922
XXB19A871F1008 5 4 23 25 40 89 79 84 nor $T=716 1514 1 0 $X=1343 $Y=922
XXB19A871F1009 5 4 26 27 42 90 79 84 nor $T=44 1514 1 0 $X=672 $Y=922
XXB19A871F1010 5 4 28 27 40 91 79 84 nor $T=-628 1514 1 0 $X=0 $Y=922
XXB19A871F1011 3 2 41 39 29 92 80 85 nand $T=-418 816 1 0 $X=0 $Y=-2
XXB19A871F1012 3 2 44 29 43 93 80 85 nand $T=254 816 1 0 $X=671 $Y=-2
XXB19A871F1013 3 2 45 39 30 94 80 85 nand $T=926 816 1 0 $X=1344 $Y=-2
XXB19A871F1014 3 2 46 30 43 95 80 85 nand $T=1598 816 1 0 $X=2016 $Y=-2
.ends 2to4_decoder_static
.subckt between_blocks 2 3 4 5 6 7 8 9 10 12 13
+	15 16 17 18 19 20 25 26 27 28 29
+	30 31 32 33 34 35 36 37 38 39 40
+	41 42 43 44 45 53
MM1 9 22 28 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1390 $Y=1777  $PIN_XY=1420,1882,1390,1777,1360,1882 $DEVICE_ID=1001
MM2 7 21 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1390 $Y=853  $PIN_XY=1420,958,1390,853,1360,958 $DEVICE_ID=1001
MM3 5 14 34 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1390 $Y=-71  $PIN_XY=1420,34,1390,-71,1360,34 $DEVICE_ID=1001
MM4 2 13 30 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1390 $Y=-974  $PIN_XY=1420,-890,1390,-974,1360,-890 $DEVICE_ID=1001
MM5 36 12 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1222 $Y=2260  $PIN_XY=1252,2176,1222,2260,1192,2176 $DEVICE_ID=1001
MM6 29 11 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1222 $Y=1357  $PIN_XY=1252,1252,1222,1357,1192,1252 $DEVICE_ID=1001
MM7 33 24 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1222 $Y=433  $PIN_XY=1252,328,1222,433,1192,328 $DEVICE_ID=1001
MM8 31 23 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1222 $Y=-491  $PIN_XY=1252,-596,1222,-491,1192,-596 $DEVICE_ID=1001
MM9 9 15 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=1798  $PIN_XY=916,1882,886,1798,856,1882 $DEVICE_ID=1001
MM10 7 15 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=874  $PIN_XY=916,958,886,874,856,958 $DEVICE_ID=1001
MM11 5 32 51 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=-50  $PIN_XY=916,34,886,-50,856,34 $DEVICE_ID=1001
MM12 2 16 49 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=-974  $PIN_XY=916,-890,886,-974,856,-890 $DEVICE_ID=1001
MM13 9 19 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=2239  $PIN_XY=748,2176,718,2239,688,2176 $DEVICE_ID=1001
MM14 22 20 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=1798  $PIN_XY=748,1882,718,1798,688,1882 $DEVICE_ID=1001
MM15 7 18 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=1336  $PIN_XY=748,1252,718,1336,688,1252 $DEVICE_ID=1001
MM16 21 17 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=874  $PIN_XY=748,958,718,874,688,958 $DEVICE_ID=1001
MM17 24 27 52 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=412  $PIN_XY=748,328,718,412,688,328 $DEVICE_ID=1001
MM18 51 16 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=-50  $PIN_XY=748,34,718,-50,688,34 $DEVICE_ID=1001
MM19 23 26 50 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=-512  $PIN_XY=748,-596,718,-512,688,-596 $DEVICE_ID=1001
MM20 49 25 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=-953  $PIN_XY=748,-890,718,-953,688,-890 $DEVICE_ID=1001
MM21 12 15 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=2260  $PIN_XY=580,2176,550,2260,520,2176 $DEVICE_ID=1001
MM22 11 15 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=1336  $PIN_XY=580,1252,550,1336,520,1252 $DEVICE_ID=1001
MM23 52 16 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=412  $PIN_XY=580,328,550,412,520,328 $DEVICE_ID=1001
MM24 50 16 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=-512  $PIN_XY=580,-596,550,-512,520,-596 $DEVICE_ID=1001
MM25 8 22 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=1777  $PIN_XY=1420,1712,1390,1777,1360,1712 $DEVICE_ID=1003
MM26 8 11 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=1437  $PIN_XY=1420,1422,1390,1437,1360,1422 $DEVICE_ID=1003
MM27 6 21 35 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=853  $PIN_XY=1420,788,1390,853,1360,788 $DEVICE_ID=1003
MM28 6 24 33 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=513  $PIN_XY=1420,498,1390,513,1360,498 $DEVICE_ID=1003
MM29 4 14 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=-71  $PIN_XY=1420,-136,1390,-71,1360,-136 $DEVICE_ID=1003
MM30 4 23 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1390 $Y=-411  $PIN_XY=1420,-426,1390,-411,1360,-426 $DEVICE_ID=1003
MM31 28 22 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=1697  $PIN_XY=1252,1712,1222,1697,1192,1712 $DEVICE_ID=1003
MM32 29 11 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=1357  $PIN_XY=1252,1422,1222,1357,1192,1422 $DEVICE_ID=1003
MM33 35 21 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=773  $PIN_XY=1252,788,1222,773,1192,788 $DEVICE_ID=1003
MM34 33 24 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=433  $PIN_XY=1252,498,1222,433,1192,498 $DEVICE_ID=1003
MM35 34 14 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=-151  $PIN_XY=1252,-136,1222,-151,1192,-136 $DEVICE_ID=1003
MM36 31 23 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1222 $Y=-491  $PIN_XY=1252,-426,1222,-491,1192,-426 $DEVICE_ID=1003
MM37 8 15 48 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=1798  $PIN_XY=916,1712,886,1798,856,1712 $DEVICE_ID=1003
MM38 6 15 46 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=874  $PIN_XY=916,788,886,874,856,788 $DEVICE_ID=1003
MM39 4 32 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=886 $Y=-50  $PIN_XY=916,-136,886,-50,856,-136 $DEVICE_ID=1003
MM40 48 20 22 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=1798  $PIN_XY=748,1712,718,1798,688,1712 $DEVICE_ID=1003
MM41 11 18 47 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=1336  $PIN_XY=748,1422,718,1336,688,1422 $DEVICE_ID=1003
MM42 46 17 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=874  $PIN_XY=748,788,718,874,688,788 $DEVICE_ID=1003
MM43 6 27 24 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=412  $PIN_XY=748,498,718,412,688,498 $DEVICE_ID=1003
MM44 14 16 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=718 $Y=-50  $PIN_XY=748,-136,718,-50,688,-136 $DEVICE_ID=1003
MM45 4 26 23 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=718 $Y=-512  $PIN_XY=748,-426,718,-512,688,-426 $DEVICE_ID=1003
MM46 47 15 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=1336  $PIN_XY=580,1422,550,1336,520,1422 $DEVICE_ID=1003
MM47 24 16 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=412  $PIN_XY=580,498,550,412,520,498 $DEVICE_ID=1003
MM48 23 16 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=550 $Y=-512  $PIN_XY=580,-426,550,-512,520,-426 $DEVICE_ID=1003
XXB19A871F1015 2 3 30 13 37 41 inv $T=1612 -680 0 180 $X=1000 $Y=-1270
XXB19A871F1016 2 4 31 23 37 42 inv $T=1000 -806 0 0 $X=1000 $Y=-806
XXB19A871F1017 5 4 34 14 38 42 inv $T=1612 244 0 180 $X=1000 $Y=-346
XXB19A871F1018 5 6 33 24 38 43 inv $T=1000 118 0 0 $X=1000 $Y=118
XXB19A871F1019 7 6 35 21 39 43 inv $T=1612 1168 0 180 $X=1000 $Y=578
XXB19A871F1020 7 8 29 11 39 44 inv $T=1000 1042 0 0 $X=1000 $Y=1042
XXB19A871F1021 9 8 28 22 40 44 inv $T=1612 2092 0 180 $X=1000 $Y=1502
XXB19A871F1022 9 10 36 12 40 45 inv $T=1000 1966 0 0 $X=1000 $Y=1966
XXB19A871F1023 7 6 21 17 15 46 39 43 nor $T=1736 1170 0 180 $X=328 $Y=578
XXB19A871F1024 7 8 11 18 15 47 39 44 nor $T=-300 1040 0 0 $X=328 $Y=1042
XXB19A871F1025 9 8 22 20 15 48 40 44 nor $T=1736 2094 0 180 $X=328 $Y=1501
XXB19A871F1026 9 10 12 19 15 53 40 45 nor $T=-300 1964 0 0 $X=328 $Y=1966
XXB19A871F1027 2 3 13 16 25 49 37 41 nand $T=1526 -452 0 180 $X=328 $Y=-1270
XXB19A871F1028 2 4 23 16 26 50 37 42 nand $T=-90 -1034 0 0 $X=327 $Y=-806
XXB19A871F1029 5 4 14 32 16 51 38 42 nand $T=1526 472 0 180 $X=328 $Y=-346
XXB19A871F1030 5 6 24 16 27 52 38 43 nand $T=-90 -110 0 0 $X=327 $Y=118
.ends between_blocks
.subckt read_circuit 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16
XXB19A871F1040 2 3 5 4 14 15 invx4 $T=-24 4 0 0 $X=0 $Y=4
XXB19A871F1041 2 3 8 7 14 15 inv $T=1512 4 0 0 $X=1512 $Y=4
XXB19A871F1042 2 3 7 5 6 16 14 15 nand $T=422 -224 0 0 $X=840 $Y=4
.ends read_circuit
.subckt buffer_highdrive 2 3 4 5 6 7 8 9
XXB19A871F1043 3 2 5 6 8 9 invx4 $T=-22 -2 0 0 $X=2 $Y=-2
XXB19A871F1044 3 2 4 5 8 9 invx4 $T=818 -2 0 0 $X=842 $Y=-2
.ends buffer_highdrive
.subckt buffer 2 3 4 5 6 7 8
XXB19A871F1045 2 3 5 4 7 8 inv $T=584 2 0 0 $X=584 $Y=2
XXB19A871F1046 2 3 4 6 7 8 inv $T=80 2 0 0 $X=80 $Y=2
.ends buffer
.subckt Demux 2 3 4 5 6 7 8 9 10 11 12
+	13 14
MM1 11 9 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1398 $Y=735  $PIN_XY=1428,672,1398,735,1368,672 $DEVICE_ID=1001
MM2 10 8 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1398 $Y=315  $PIN_XY=1428,378,1398,315,1368,378 $DEVICE_ID=1001
MM3 9 6 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=894 $Y=735  $PIN_XY=924,672,894,735,864,672 $DEVICE_ID=1001
MM4 8 5 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=894 $Y=315  $PIN_XY=924,378,894,315,864,378 $DEVICE_ID=1001
MM5 15 7 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=726 $Y=735  $PIN_XY=756,672,726,735,696,672 $DEVICE_ID=1001
MM6 16 7 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=726 $Y=315  $PIN_XY=756,378,726,315,696,378 $DEVICE_ID=1001
MM7 6 5 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=756  $PIN_XY=252,672,222,756,192,672 $DEVICE_ID=1001
XXB19A871F1047 2 3 _GENERATED_17 2 12 13 sram_filler $T=616 588 0 180 $X=167 $Y=-2
XXB19A871F1048 2 3 3 _GENERATED_18 12 13 sram_filler $T=448 588 0 180 $X=0 $Y=-2
XXB19A871F1049 2 4 6 5 12 14 inv $T=0 462 0 0 $X=0 $Y=462
XXB19A871F1050 2 4 11 9 12 14 inv $T=1176 462 0 0 $X=1176 $Y=462
XXB19A871F1051 2 3 10 8 12 13 inv $T=1176 588 1 0 $X=1176 $Y=-2
XXB19A871F1052 2 4 9 7 6 15 12 14 nand $T=86 234 0 0 $X=504 $Y=462
XXB19A871F1053 2 3 8 7 5 16 12 13 nand $T=86 816 1 0 $X=504 $Y=-2
.ends Demux

* Hierarchy Level 1
.subckt static_row_decoder_3by8 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16 17 18 26 27 28 31 32
+	34 51 52 53 54 55 56 57 58 59 60
+	61 62 63 64 65 66 67 68 69 70 71
+	72 73 74 75 88 112
*.floating_nets 107 108 109 110 111
MM1 16 90 57 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=884  $PIN_XY=3760,800,3730,884,3700,800 $DEVICE_ID=1001
MM2 11 91 58 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-40  $PIN_XY=3760,-124,3730,-40,3700,-124 $DEVICE_ID=1001
MM3 10 87 54 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-964  $PIN_XY=3760,-1048,3730,-964,3700,-1048 $DEVICE_ID=1001
MM4 13 86 53 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-1888  $PIN_XY=3760,-1972,3730,-1888,3700,-1972 $DEVICE_ID=1001
MM5 5 84 51 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-2812  $PIN_XY=3760,-2896,3730,-2812,3700,-2896 $DEVICE_ID=1001
MM6 8 89 56 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-3736  $PIN_XY=3760,-3820,3730,-3736,3700,-3820 $DEVICE_ID=1001
MM7 3 85 52 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3730 $Y=-4660  $PIN_XY=3760,-4744,3730,-4660,3700,-4744 $DEVICE_ID=1001
MM8 57 90 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=884  $PIN_XY=3592,800,3562,884,3532,800 $DEVICE_ID=1001
MM9 58 91 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-40  $PIN_XY=3592,-124,3562,-40,3532,-124 $DEVICE_ID=1001
MM10 54 87 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-964  $PIN_XY=3592,-1048,3562,-964,3532,-1048 $DEVICE_ID=1001
MM11 53 86 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-1888  $PIN_XY=3592,-1972,3562,-1888,3532,-1972 $DEVICE_ID=1001
MM12 51 84 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-2812  $PIN_XY=3592,-2896,3562,-2812,3532,-2896 $DEVICE_ID=1001
MM13 56 89 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-3736  $PIN_XY=3592,-3820,3562,-3736,3532,-3820 $DEVICE_ID=1001
MM14 52 85 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-4660  $PIN_XY=3592,-4744,3562,-4660,3532,-4744 $DEVICE_ID=1001
MM15 15 50 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=1346  $PIN_XY=2920,1430,2890,1346,2860,1430 $DEVICE_ID=1001
MM16 16 25 90 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=884  $PIN_XY=2920,800,2890,884,2860,800 $DEVICE_ID=1001
MM17 16 49 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=422  $PIN_XY=2920,506,2890,422,2860,506 $DEVICE_ID=1001
MM18 11 24 91 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-40  $PIN_XY=2920,-124,2890,-40,2860,-124 $DEVICE_ID=1001
MM19 11 48 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-502  $PIN_XY=2920,-418,2890,-502,2860,-418 $DEVICE_ID=1001
MM20 10 23 87 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-964  $PIN_XY=2920,-1048,2890,-964,2860,-1048 $DEVICE_ID=1001
MM21 10 47 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-1426  $PIN_XY=2920,-1342,2890,-1426,2860,-1342 $DEVICE_ID=1001
MM22 13 22 86 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-1888  $PIN_XY=2920,-1972,2890,-1888,2860,-1972 $DEVICE_ID=1001
MM23 13 43 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-2350  $PIN_XY=2920,-2266,2890,-2350,2860,-2266 $DEVICE_ID=1001
MM24 5 21 84 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-2812  $PIN_XY=2920,-2896,2890,-2812,2860,-2896 $DEVICE_ID=1001
MM25 5 42 20 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-3274  $PIN_XY=2920,-3190,2890,-3274,2860,-3190 $DEVICE_ID=1001
MM26 8 20 89 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-3736  $PIN_XY=2920,-3820,2890,-3736,2860,-3820 $DEVICE_ID=1001
MM27 8 41 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-4198  $PIN_XY=2920,-4114,2890,-4198,2860,-4114 $DEVICE_ID=1001
MM28 3 19 85 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-4660  $PIN_XY=2920,-4744,2890,-4660,2860,-4744 $DEVICE_ID=1001
MM29 25 46 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=1346  $PIN_XY=2752,1430,2722,1346,2692,1430 $DEVICE_ID=1001
MM30 90 25 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=884  $PIN_XY=2752,800,2722,884,2692,800 $DEVICE_ID=1001
MM31 24 45 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=422  $PIN_XY=2752,506,2722,422,2692,506 $DEVICE_ID=1001
MM32 91 24 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-40  $PIN_XY=2752,-124,2722,-40,2692,-124 $DEVICE_ID=1001
MM33 23 44 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-502  $PIN_XY=2752,-418,2722,-502,2692,-418 $DEVICE_ID=1001
MM34 87 23 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-964  $PIN_XY=2752,-1048,2722,-964,2692,-1048 $DEVICE_ID=1001
MM35 22 40 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-1426  $PIN_XY=2752,-1342,2722,-1426,2692,-1342 $DEVICE_ID=1001
MM36 86 22 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-1888  $PIN_XY=2752,-1972,2722,-1888,2692,-1972 $DEVICE_ID=1001
MM37 21 39 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-2350  $PIN_XY=2752,-2266,2722,-2350,2692,-2266 $DEVICE_ID=1001
MM38 84 21 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-2812  $PIN_XY=2752,-2896,2722,-2812,2692,-2896 $DEVICE_ID=1001
MM39 20 38 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-3274  $PIN_XY=2752,-3190,2722,-3274,2692,-3190 $DEVICE_ID=1001
MM40 89 20 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-3736  $PIN_XY=2752,-3820,2722,-3736,2692,-3820 $DEVICE_ID=1001
MM41 19 37 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-4198  $PIN_XY=2752,-4114,2722,-4198,2692,-4114 $DEVICE_ID=1001
MM42 85 19 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-4660  $PIN_XY=2752,-4744,2722,-4660,2692,-4744 $DEVICE_ID=1001
MM43 50 36 105 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=1346  $PIN_XY=2248,1430,2218,1346,2188,1430 $DEVICE_ID=1001
MM44 46 28 106 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=884  $PIN_XY=2248,800,2218,884,2188,800 $DEVICE_ID=1001
MM45 49 36 104 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=422  $PIN_XY=2248,506,2218,422,2188,506 $DEVICE_ID=1001
MM46 45 28 99 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-40  $PIN_XY=2248,-124,2218,-40,2188,-124 $DEVICE_ID=1001
MM47 48 27 102 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-502  $PIN_XY=2248,-418,2218,-502,2188,-418 $DEVICE_ID=1001
MM48 44 28 103 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-964  $PIN_XY=2248,-1048,2218,-964,2188,-1048 $DEVICE_ID=1001
MM49 47 27 101 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-1426  $PIN_XY=2248,-1342,2218,-1426,2188,-1342 $DEVICE_ID=1001
MM50 40 28 100 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-1888  $PIN_XY=2248,-1972,2218,-1888,2188,-1972 $DEVICE_ID=1001
MM51 43 36 93 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-2350  $PIN_XY=2248,-2266,2218,-2350,2188,-2266 $DEVICE_ID=1001
MM52 39 28 92 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-2812  $PIN_XY=2248,-2896,2218,-2812,2188,-2896 $DEVICE_ID=1001
MM53 42 36 94 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-3274  $PIN_XY=2248,-3190,2218,-3274,2188,-3190 $DEVICE_ID=1001
MM54 38 28 95 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-3736  $PIN_XY=2248,-3820,2218,-3736,2188,-3820 $DEVICE_ID=1001
MM55 41 27 97 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-4198  $PIN_XY=2248,-4114,2218,-4198,2188,-4114 $DEVICE_ID=1001
MM56 37 28 96 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-4660  $PIN_XY=2248,-4744,2218,-4660,2188,-4744 $DEVICE_ID=1001
MM57 105 29 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=1346  $PIN_XY=2080,1430,2050,1346,2020,1430 $DEVICE_ID=1001
MM58 106 35 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=884  $PIN_XY=2080,800,2050,884,2020,800 $DEVICE_ID=1001
MM59 104 26 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=422  $PIN_XY=2080,506,2050,422,2020,506 $DEVICE_ID=1001
MM60 99 35 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-40  $PIN_XY=2080,-124,2050,-40,2020,-124 $DEVICE_ID=1001
MM61 102 29 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-502  $PIN_XY=2080,-418,2050,-502,2020,-418 $DEVICE_ID=1001
MM62 103 35 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-964  $PIN_XY=2080,-1048,2050,-964,2020,-1048 $DEVICE_ID=1001
MM63 101 26 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-1426  $PIN_XY=2080,-1342,2050,-1426,2020,-1342 $DEVICE_ID=1001
MM64 100 35 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-1888  $PIN_XY=2080,-1972,2050,-1888,2020,-1972 $DEVICE_ID=1001
MM65 93 29 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-2350  $PIN_XY=2080,-2266,2050,-2350,2020,-2266 $DEVICE_ID=1001
MM66 92 31 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-2812  $PIN_XY=2080,-2896,2050,-2812,2020,-2896 $DEVICE_ID=1001
MM67 94 31 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-3274  $PIN_XY=2080,-3190,2050,-3274,2020,-3190 $DEVICE_ID=1001
MM68 95 26 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-3736  $PIN_XY=2080,-3820,2050,-3736,2020,-3820 $DEVICE_ID=1001
MM69 97 29 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-4198  $PIN_XY=2080,-4114,2050,-4198,2020,-4114 $DEVICE_ID=1001
MM70 96 31 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-4660  $PIN_XY=2080,-4744,2050,-4660,2020,-4744 $DEVICE_ID=1001
MM71 29 26 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1546 $Y=1346  $PIN_XY=1576,1430,1546,1346,1516,1430 $DEVICE_ID=1001
MM72 36 27 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1546 $Y=884  $PIN_XY=1576,800,1546,884,1516,800 $DEVICE_ID=1001
MM73 35 31 16 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1546 $Y=443  $PIN_XY=1576,506,1546,443,1516,506 $DEVICE_ID=1001
MM74 3 34 30 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1042 $Y=-4681  $PIN_XY=1072,-4744,1042,-4681,1012,-4744 $DEVICE_ID=1001
MM75 30 34 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=874 $Y=-4681  $PIN_XY=904,-4744,874,-4681,844,-4744 $DEVICE_ID=1001
MM76 3 33 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-5122  $PIN_XY=2920,-5038,2890,-5122,2860,-5038 $DEVICE_ID=1001
MM77 18 32 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-5122  $PIN_XY=2752,-5038,2722,-5122,2692,-5038 $DEVICE_ID=1001
MM78 33 27 98 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-5122  $PIN_XY=2248,-5038,2218,-5122,2188,-5038 $DEVICE_ID=1001
MM79 98 31 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-5122  $PIN_XY=2080,-5038,2050,-5122,2020,-5038 $DEVICE_ID=1001
MM80 3 30 28 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1042 $Y=-5101  $PIN_XY=1072,-5038,1042,-5101,1012,-5038 $DEVICE_ID=1001
MM81 28 30 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=874 $Y=-5101  $PIN_XY=904,-5038,874,-5101,844,-5038 $DEVICE_ID=1001
MM82 14 90 57 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=964  $PIN_XY=4096,970,4066,964,4036,970 $DEVICE_ID=1003
MM83 17 91 58 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=40  $PIN_XY=4096,46,4066,40,4036,46 $DEVICE_ID=1003
MM84 9 87 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-884  $PIN_XY=4096,-878,4066,-884,4036,-878 $DEVICE_ID=1003
MM85 12 86 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-1808  $PIN_XY=4096,-1802,4066,-1808,4036,-1802 $DEVICE_ID=1003
MM86 6 84 51 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-2732  $PIN_XY=4096,-2726,4066,-2732,4036,-2726 $DEVICE_ID=1003
MM87 7 89 56 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-3656  $PIN_XY=4096,-3650,4066,-3656,4036,-3650 $DEVICE_ID=1003
MM88 2 85 52 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-4580  $PIN_XY=4096,-4574,4066,-4580,4036,-4574 $DEVICE_ID=1003
MM89 57 90 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=964  $PIN_XY=3928,970,3898,964,3868,970 $DEVICE_ID=1003
MM90 58 91 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=40  $PIN_XY=3928,46,3898,40,3868,46 $DEVICE_ID=1003
MM91 54 87 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-884  $PIN_XY=3928,-878,3898,-884,3868,-878 $DEVICE_ID=1003
MM92 53 86 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-1808  $PIN_XY=3928,-1802,3898,-1808,3868,-1802 $DEVICE_ID=1003
MM93 51 84 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-2732  $PIN_XY=3928,-2726,3898,-2732,3868,-2726 $DEVICE_ID=1003
MM94 56 89 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-3656  $PIN_XY=3928,-3650,3898,-3656,3868,-3650 $DEVICE_ID=1003
MM95 52 85 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-4580  $PIN_XY=3928,-4574,3898,-4580,3868,-4574 $DEVICE_ID=1003
MM96 14 90 57 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=884  $PIN_XY=3760,970,3730,884,3700,970 $DEVICE_ID=1003
MM97 17 91 58 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-40  $PIN_XY=3760,46,3730,-40,3700,46 $DEVICE_ID=1003
MM98 9 87 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-964  $PIN_XY=3760,-878,3730,-964,3700,-878 $DEVICE_ID=1003
MM99 12 86 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-1888  $PIN_XY=3760,-1802,3730,-1888,3700,-1802 $DEVICE_ID=1003
MM100 6 84 51 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-2812  $PIN_XY=3760,-2726,3730,-2812,3700,-2726 $DEVICE_ID=1003
MM101 7 89 56 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-3736  $PIN_XY=3760,-3650,3730,-3736,3700,-3650 $DEVICE_ID=1003
MM102 57 90 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=884  $PIN_XY=3592,970,3562,884,3532,970 $DEVICE_ID=1003
MM103 58 91 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-40  $PIN_XY=3592,46,3562,-40,3532,46 $DEVICE_ID=1003
MM104 54 87 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-964  $PIN_XY=3592,-878,3562,-964,3532,-878 $DEVICE_ID=1003
MM105 53 86 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-1888  $PIN_XY=3592,-1802,3562,-1888,3532,-1802 $DEVICE_ID=1003
MM106 51 84 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-2812  $PIN_XY=3592,-2726,3562,-2812,3532,-2726 $DEVICE_ID=1003
MM107 56 89 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-3736  $PIN_XY=3592,-3650,3562,-3736,3532,-3650 $DEVICE_ID=1003
MM108 14 25 90 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=964  $PIN_XY=3256,970,3226,964,3196,970 $DEVICE_ID=1003
MM109 17 24 91 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=40  $PIN_XY=3256,46,3226,40,3196,46 $DEVICE_ID=1003
MM110 9 23 87 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-884  $PIN_XY=3256,-878,3226,-884,3196,-878 $DEVICE_ID=1003
MM111 12 22 86 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-1808  $PIN_XY=3256,-1802,3226,-1808,3196,-1802 $DEVICE_ID=1003
MM112 6 21 84 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-2732  $PIN_XY=3256,-2726,3226,-2732,3196,-2726 $DEVICE_ID=1003
MM113 7 20 89 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-3656  $PIN_XY=3256,-3650,3226,-3656,3196,-3650 $DEVICE_ID=1003
MM114 2 19 85 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-4580  $PIN_XY=3256,-4574,3226,-4580,3196,-4574 $DEVICE_ID=1003
MM115 90 25 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=964  $PIN_XY=3088,970,3058,964,3028,970 $DEVICE_ID=1003
MM116 91 24 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=40  $PIN_XY=3088,46,3058,40,3028,46 $DEVICE_ID=1003
MM117 87 23 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-884  $PIN_XY=3088,-878,3058,-884,3028,-878 $DEVICE_ID=1003
MM118 86 22 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-1808  $PIN_XY=3088,-1802,3058,-1808,3028,-1802 $DEVICE_ID=1003
MM119 84 21 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-2732  $PIN_XY=3088,-2726,3058,-2732,3028,-2726 $DEVICE_ID=1003
MM120 89 20 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-3656  $PIN_XY=3088,-3650,3058,-3656,3028,-3650 $DEVICE_ID=1003
MM121 85 19 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-4580  $PIN_XY=3088,-4574,3058,-4580,3028,-4574 $DEVICE_ID=1003
MM122 25 50 82 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=1346  $PIN_XY=2920,1260,2890,1346,2860,1260 $DEVICE_ID=1003
MM123 14 25 90 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=884  $PIN_XY=2920,970,2890,884,2860,970 $DEVICE_ID=1003
MM124 24 49 83 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=422  $PIN_XY=2920,336,2890,422,2860,336 $DEVICE_ID=1003
MM125 17 24 91 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-40  $PIN_XY=2920,46,2890,-40,2860,46 $DEVICE_ID=1003
MM126 23 48 81 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-502  $PIN_XY=2920,-588,2890,-502,2860,-588 $DEVICE_ID=1003
MM127 9 23 87 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-964  $PIN_XY=2920,-878,2890,-964,2860,-878 $DEVICE_ID=1003
MM128 22 47 80 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-1426  $PIN_XY=2920,-1512,2890,-1426,2860,-1512 $DEVICE_ID=1003
MM129 12 22 86 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-1888  $PIN_XY=2920,-1802,2890,-1888,2860,-1802 $DEVICE_ID=1003
MM130 21 43 77 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-2350  $PIN_XY=2920,-2436,2890,-2350,2860,-2436 $DEVICE_ID=1003
MM131 6 21 84 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-2812  $PIN_XY=2920,-2726,2890,-2812,2860,-2726 $DEVICE_ID=1003
MM132 20 42 78 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-3274  $PIN_XY=2920,-3360,2890,-3274,2860,-3360 $DEVICE_ID=1003
MM133 7 20 89 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-3736  $PIN_XY=2920,-3650,2890,-3736,2860,-3650 $DEVICE_ID=1003
MM134 19 41 76 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-4198  $PIN_XY=2920,-4284,2890,-4198,2860,-4284 $DEVICE_ID=1003
MM135 82 46 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=1346  $PIN_XY=2752,1260,2722,1346,2692,1260 $DEVICE_ID=1003
MM136 90 25 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=884  $PIN_XY=2752,970,2722,884,2692,970 $DEVICE_ID=1003
MM137 83 45 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=422  $PIN_XY=2752,336,2722,422,2692,336 $DEVICE_ID=1003
MM138 91 24 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-40  $PIN_XY=2752,46,2722,-40,2692,46 $DEVICE_ID=1003
MM139 81 44 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-502  $PIN_XY=2752,-588,2722,-502,2692,-588 $DEVICE_ID=1003
MM140 87 23 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-964  $PIN_XY=2752,-878,2722,-964,2692,-878 $DEVICE_ID=1003
MM141 80 40 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-1426  $PIN_XY=2752,-1512,2722,-1426,2692,-1512 $DEVICE_ID=1003
MM142 86 22 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-1888  $PIN_XY=2752,-1802,2722,-1888,2692,-1802 $DEVICE_ID=1003
MM143 77 39 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-2350  $PIN_XY=2752,-2436,2722,-2350,2692,-2436 $DEVICE_ID=1003
MM144 84 21 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-2812  $PIN_XY=2752,-2726,2722,-2812,2692,-2726 $DEVICE_ID=1003
MM145 78 38 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-3274  $PIN_XY=2752,-3360,2722,-3274,2692,-3360 $DEVICE_ID=1003
MM146 89 20 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-3736  $PIN_XY=2752,-3650,2722,-3736,2692,-3650 $DEVICE_ID=1003
MM147 76 37 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-4198  $PIN_XY=2752,-4284,2722,-4198,2692,-4284 $DEVICE_ID=1003
MM148 14 36 50 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=1346  $PIN_XY=2248,1260,2218,1346,2188,1260 $DEVICE_ID=1003
MM149 14 28 46 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=884  $PIN_XY=2248,970,2218,884,2188,970 $DEVICE_ID=1003
MM150 17 36 49 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=422  $PIN_XY=2248,336,2218,422,2188,336 $DEVICE_ID=1003
MM151 17 28 45 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-40  $PIN_XY=2248,46,2218,-40,2188,46 $DEVICE_ID=1003
MM152 9 27 48 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-502  $PIN_XY=2248,-588,2218,-502,2188,-588 $DEVICE_ID=1003
MM153 9 28 44 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-964  $PIN_XY=2248,-878,2218,-964,2188,-878 $DEVICE_ID=1003
MM154 12 27 47 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-1426  $PIN_XY=2248,-1512,2218,-1426,2188,-1512 $DEVICE_ID=1003
MM155 12 28 40 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-1888  $PIN_XY=2248,-1802,2218,-1888,2188,-1802 $DEVICE_ID=1003
MM156 6 36 43 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-2350  $PIN_XY=2248,-2436,2218,-2350,2188,-2436 $DEVICE_ID=1003
MM157 6 28 39 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-2812  $PIN_XY=2248,-2726,2218,-2812,2188,-2726 $DEVICE_ID=1003
MM158 7 36 42 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-3274  $PIN_XY=2248,-3360,2218,-3274,2188,-3360 $DEVICE_ID=1003
MM159 7 28 38 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-3736  $PIN_XY=2248,-3650,2218,-3736,2188,-3650 $DEVICE_ID=1003
MM160 2 27 41 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-4198  $PIN_XY=2248,-4284,2218,-4198,2188,-4284 $DEVICE_ID=1003
MM161 50 29 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=1346  $PIN_XY=2080,1260,2050,1346,2020,1260 $DEVICE_ID=1003
MM162 46 35 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=884  $PIN_XY=2080,970,2050,884,2020,970 $DEVICE_ID=1003
MM163 49 26 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=422  $PIN_XY=2080,336,2050,422,2020,336 $DEVICE_ID=1003
MM164 45 35 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-40  $PIN_XY=2080,46,2050,-40,2020,46 $DEVICE_ID=1003
MM165 48 29 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-502  $PIN_XY=2080,-588,2050,-502,2020,-588 $DEVICE_ID=1003
MM166 44 35 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-964  $PIN_XY=2080,-878,2050,-964,2020,-878 $DEVICE_ID=1003
MM167 47 26 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-1426  $PIN_XY=2080,-1512,2050,-1426,2020,-1512 $DEVICE_ID=1003
MM168 40 35 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-1888  $PIN_XY=2080,-1802,2050,-1888,2020,-1802 $DEVICE_ID=1003
MM169 43 29 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-2350  $PIN_XY=2080,-2436,2050,-2350,2020,-2436 $DEVICE_ID=1003
MM170 39 31 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-2812  $PIN_XY=2080,-2726,2050,-2812,2020,-2726 $DEVICE_ID=1003
MM171 42 31 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-3274  $PIN_XY=2080,-3360,2050,-3274,2020,-3360 $DEVICE_ID=1003
MM172 38 26 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-3736  $PIN_XY=2080,-3650,2050,-3736,2020,-3650 $DEVICE_ID=1003
MM173 41 29 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-4198  $PIN_XY=2080,-4284,2050,-4198,2020,-4284 $DEVICE_ID=1003
MM174 14 26 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1714 $Y=1245  $PIN_XY=1744,1260,1714,1245,1684,1260 $DEVICE_ID=1003
MM175 14 27 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1714 $Y=985  $PIN_XY=1744,970,1714,985,1684,970 $DEVICE_ID=1003
MM176 17 31 35 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1714 $Y=342  $PIN_XY=1744,336,1714,342,1684,336 $DEVICE_ID=1003
MM177 29 26 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1546 $Y=1346  $PIN_XY=1576,1260,1546,1346,1516,1260 $DEVICE_ID=1003
MM178 36 27 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1546 $Y=884  $PIN_XY=1576,970,1546,884,1516,970 $DEVICE_ID=1003
MM179 35 31 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1546 $Y=443  $PIN_XY=1576,336,1546,443,1516,336 $DEVICE_ID=1003
MM180 2 34 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1378 $Y=-4580  $PIN_XY=1408,-4574,1378,-4580,1348,-4574 $DEVICE_ID=1003
MM181 30 34 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1210 $Y=-4580  $PIN_XY=1240,-4574,1210,-4580,1180,-4574 $DEVICE_ID=1003
MM182 2 88 55 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4066 $Y=-5504  $PIN_XY=4096,-5498,4066,-5504,4036,-5498 $DEVICE_ID=1003
MM183 55 88 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3898 $Y=-5504  $PIN_XY=3928,-5498,3898,-5504,3868,-5498 $DEVICE_ID=1003
MM184 2 85 52 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-4660  $PIN_XY=3760,-4574,3730,-4660,3700,-4574 $DEVICE_ID=1003
MM185 2 88 55 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3730 $Y=-5584  $PIN_XY=3760,-5498,3730,-5584,3700,-5498 $DEVICE_ID=1003
MM186 52 85 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-4660  $PIN_XY=3592,-4574,3562,-4660,3532,-4574 $DEVICE_ID=1003
MM187 55 88 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3562 $Y=-5584  $PIN_XY=3592,-5498,3562,-5584,3532,-5498 $DEVICE_ID=1003
MM188 2 18 88 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3226 $Y=-5504  $PIN_XY=3256,-5498,3226,-5504,3196,-5498 $DEVICE_ID=1003
MM189 88 18 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3058 $Y=-5504  $PIN_XY=3088,-5498,3058,-5504,3028,-5498 $DEVICE_ID=1003
MM190 2 19 85 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-4660  $PIN_XY=2920,-4574,2890,-4660,2860,-4574 $DEVICE_ID=1003
MM191 18 33 79 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2890 $Y=-5122  $PIN_XY=2920,-5208,2890,-5122,2860,-5208 $DEVICE_ID=1003
MM192 2 18 88 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2890 $Y=-5563  $PIN_XY=2920,-5498,2890,-5563,2860,-5498 $DEVICE_ID=1003
MM193 85 19 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-4660  $PIN_XY=2752,-4574,2722,-4660,2692,-4574 $DEVICE_ID=1003
MM194 79 32 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-5122  $PIN_XY=2752,-5208,2722,-5122,2692,-5208 $DEVICE_ID=1003
MM195 88 18 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2722 $Y=-5563  $PIN_XY=2752,-5498,2722,-5563,2692,-5498 $DEVICE_ID=1003
MM196 2 28 37 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-4660  $PIN_XY=2248,-4574,2218,-4660,2188,-4574 $DEVICE_ID=1003
MM197 2 27 33 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-5122  $PIN_XY=2248,-5208,2218,-5122,2188,-5208 $DEVICE_ID=1003
MM198 2 28 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2218 $Y=-5563  $PIN_XY=2248,-5498,2218,-5563,2188,-5498 $DEVICE_ID=1003
MM199 37 31 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-4660  $PIN_XY=2080,-4574,2050,-4660,2020,-4574 $DEVICE_ID=1003
MM200 33 31 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-5122  $PIN_XY=2080,-5208,2050,-5122,2020,-5208 $DEVICE_ID=1003
MM201 32 26 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2050 $Y=-5563  $PIN_XY=2080,-5498,2050,-5563,2020,-5498 $DEVICE_ID=1003
MM202 2 30 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1378 $Y=-5202  $PIN_XY=1408,-5208,1378,-5202,1348,-5208 $DEVICE_ID=1003
MM203 28 30 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1210 $Y=-5202  $PIN_XY=1240,-5208,1210,-5202,1180,-5208 $DEVICE_ID=1003
MM204 2 34 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1042 $Y=-4681  $PIN_XY=1072,-4574,1042,-4681,1012,-4574 $DEVICE_ID=1003
MM205 2 30 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1042 $Y=-5101  $PIN_XY=1072,-5208,1042,-5101,1012,-5208 $DEVICE_ID=1003
MM206 30 34 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=874 $Y=-4681  $PIN_XY=904,-4574,874,-4681,844,-4574 $DEVICE_ID=1003
MM207 28 30 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=874 $Y=-5101  $PIN_XY=904,-5208,874,-5101,844,-5208 $DEVICE_ID=1003
XXB19A871F772 16 17 35 31 66 73 inv $T=1324 716 1 0 $X=1324 $Y=126
XXB19A871F773 15 14 29 26 65 75 inv $T=1324 1640 1 0 $X=1324 $Y=1050
XXB19A871F774 16 14 36 27 66 75 inv $T=1324 590 0 0 $X=1324 $Y=590
XXB19A871F775 8 2 19 41 37 76 62 69 nor $T=1872 -3902 1 0 $X=2500 $Y=-4494
XXB19A871F776 13 6 21 43 39 77 64 71 nor $T=1872 -2054 1 0 $X=2500 $Y=-2646
XXB19A871F777 5 7 20 42 38 78 61 70 nor $T=1872 -2978 1 0 $X=2500 $Y=-3570
XXB19A871F778 3 2 18 33 32 79 60 68 nor $T=1872 -4826 1 0 $X=2500 $Y=-5418
XXB19A871F779 10 12 22 47 40 80 63 72 nor $T=1872 -1130 1 0 $X=2500 $Y=-1722
XXB19A871F780 11 9 23 48 44 81 67 74 nor $T=1872 -206 1 0 $X=2500 $Y=-798
XXB19A871F781 15 14 25 50 46 82 65 75 nor $T=1872 1642 1 0 $X=2500 $Y=1050
XXB19A871F782 16 17 24 49 45 83 66 73 nor $T=1872 718 1 0 $X=2500 $Y=126
XXB19A871F783 5 6 39 31 28 92 61 71 nand $T=1410 -3334 0 0 $X=1827 $Y=-3106
XXB19A871F784 13 6 43 29 36 93 64 71 nand $T=1410 -1828 1 0 $X=1827 $Y=-2646
XXB19A871F785 5 7 42 31 36 94 61 70 nand $T=1410 -2752 1 0 $X=1827 $Y=-3570
XXB19A871F786 8 7 38 26 28 95 62 70 nand $T=1410 -4258 0 0 $X=1827 $Y=-4030
XXB19A871F787 4 2 32 26 28 112 59 68 nand $T=1410 -6106 0 0 $X=1827 $Y=-5878
XXB19A871F788 3 2 37 31 28 96 60 69 nand $T=1410 -5182 0 0 $X=1827 $Y=-4954
XXB19A871F789 8 2 41 29 27 97 62 69 nand $T=1410 -3676 1 0 $X=1827 $Y=-4494
XXB19A871F790 3 2 33 31 27 98 60 68 nand $T=1410 -4600 1 0 $X=1827 $Y=-5418
XXB19A871F791 11 17 45 35 28 99 67 73 nand $T=1410 -562 0 0 $X=1827 $Y=-334
XXB19A871F792 13 12 40 35 28 100 64 72 nand $T=1410 -2410 0 0 $X=1827 $Y=-2182
XXB19A871F793 10 12 47 26 27 101 63 72 nand $T=1410 -904 1 0 $X=1827 $Y=-1722
XXB19A871F794 11 9 48 29 27 102 67 74 nand $T=1410 20 1 0 $X=1827 $Y=-798
XXB19A871F795 10 9 44 35 28 103 63 74 nand $T=1410 -1486 0 0 $X=1827 $Y=-1258
XXB19A871F796 16 17 49 26 36 104 66 73 nand $T=1410 944 1 0 $X=1827 $Y=126
XXB19A871F797 15 14 50 29 36 105 65 75 nand $T=1410 1868 1 0 $X=1827 $Y=1050
XXB19A871F798 16 14 46 35 28 106 66 75 nand $T=1410 362 0 0 $X=1827 $Y=590
XXB19A871F799 6 5 51 84 21 39 61 71 buffer_highdrive $T=2498 -3104 0 0 $X=2500 $Y=-3106
XXB19A871F800 2 3 52 85 19 37 60 69 buffer_highdrive $T=2498 -4952 0 0 $X=2500 $Y=-4954
XXB19A871F801 12 13 53 86 22 40 64 72 buffer_highdrive $T=2498 -2180 0 0 $X=2500 $Y=-2182
XXB19A871F802 9 10 54 87 23 44 63 74 buffer_highdrive $T=2498 -1256 0 0 $X=2500 $Y=-1258
XXB19A871F803 2 4 55 88 18 32 59 68 buffer_highdrive $T=2498 -5876 0 0 $X=2500 $Y=-5878
XXB19A871F804 7 8 56 89 20 38 62 70 buffer_highdrive $T=2498 -4028 0 0 $X=2500 $Y=-4030
XXB19A871F805 14 16 57 90 25 46 66 75 buffer_highdrive $T=2498 592 0 0 $X=2500 $Y=590
XXB19A871F806 17 11 58 91 24 45 67 73 buffer_highdrive $T=2498 -332 0 0 $X=2500 $Y=-334
XXB19A871F807 3 2 28 30 60 68 invx4 $T=628 -4828 1 0 $X=652 $Y=-5418
XXB19A871F808 3 2 30 34 60 69 invx4 $T=628 -4954 0 0 $X=652 $Y=-4954
XXB19A871F809 15 14 _GENERATED_114 _GENERATED_113 65 75 sram_filler $T=1100 1640 0 180 $X=652 $Y=1050
XXB19A871F810 16 14 _GENERATED_116 _GENERATED_115 66 75 sram_filler $T=648 590 0 0 $X=652 $Y=590
XXB19A871F811 16 17 _GENERATED_118 _GENERATED_117 66 73 sram_filler $T=1100 716 0 180 $X=652 $Y=126
XXB19A871F812 16 17 _GENERATED_120 _GENERATED_119 66 73 sram_filler $T=1436 716 0 180 $X=988 $Y=126
XXB19A871F813 16 14 _GENERATED_122 _GENERATED_121 66 75 sram_filler $T=984 590 0 0 $X=988 $Y=590
XXB19A871F814 15 14 _GENERATED_124 _GENERATED_123 65 75 sram_filler $T=1436 1640 0 180 $X=988 $Y=1050
XXB19A871F815 4 2 _GENERATED_126 _GENERATED_125 59 68 sram_filler $T=648 -5878 0 0 $X=652 $Y=-5878
XXB19A871F816 4 2 _GENERATED_128 _GENERATED_127 59 68 sram_filler $T=984 -5878 0 0 $X=988 $Y=-5878
XXB19A871F817 4 2 _GENERATED_129 4 59 68 sram_filler $T=1320 -5878 0 0 $X=1324 $Y=-5878
XXB19A871F818 4 2 2 _GENERATED_130 59 68 sram_filler $T=1488 -5878 0 0 $X=1492 $Y=-5878
XXB19A871F819 11 17 _GENERATED_132 _GENERATED_131 67 73 sram_filler $T=648 -334 0 0 $X=652 $Y=-334
XXB19A871F820 11 17 _GENERATED_134 _GENERATED_133 67 73 sram_filler $T=984 -334 0 0 $X=988 $Y=-334
XXB19A871F821 11 17 _GENERATED_135 11 67 73 sram_filler $T=1320 -334 0 0 $X=1324 $Y=-334
XXB19A871F822 11 17 17 _GENERATED_136 67 73 sram_filler $T=1488 -334 0 0 $X=1492 $Y=-334
XXB19A871F823 10 9 _GENERATED_137 10 63 74 sram_filler $T=648 -1258 0 0 $X=652 $Y=-1258
XXB19A871F824 10 9 9 _GENERATED_138 63 74 sram_filler $T=816 -1258 0 0 $X=820 $Y=-1258
XXB19A871F825 10 9 _GENERATED_140 _GENERATED_139 63 74 sram_filler $T=1152 -1258 0 0 $X=1156 $Y=-1258
XXB19A871F826 10 9 _GENERATED_142 _GENERATED_141 63 74 sram_filler $T=1488 -1258 0 0 $X=1492 $Y=-1258
XXB19A871F827 11 9 9 _GENERATED_143 67 74 sram_filler $T=1100 -208 0 180 $X=652 $Y=-798
XXB19A871F828 11 9 _GENERATED_144 11 67 74 sram_filler $T=1268 -208 0 180 $X=820 $Y=-798
XXB19A871F829 11 9 _GENERATED_146 _GENERATED_145 67 74 sram_filler $T=1604 -208 0 180 $X=1156 $Y=-798
XXB19A871F830 11 9 _GENERATED_148 _GENERATED_147 67 74 sram_filler $T=1940 -208 0 180 $X=1492 $Y=-798
XXB19A871F831 10 12 _GENERATED_150 _GENERATED_149 63 72 sram_filler $T=1940 -1132 0 180 $X=1492 $Y=-1722
XXB19A871F832 10 12 _GENERATED_152 _GENERATED_151 63 72 sram_filler $T=1604 -1132 0 180 $X=1156 $Y=-1722
XXB19A871F833 10 12 _GENERATED_153 10 63 72 sram_filler $T=1268 -1132 0 180 $X=820 $Y=-1722
XXB19A871F834 10 12 12 _GENERATED_154 63 72 sram_filler $T=1100 -1132 0 180 $X=652 $Y=-1722
XXB19A871F835 13 12 _GENERATED_156 _GENERATED_155 64 72 sram_filler $T=1488 -2182 0 0 $X=1492 $Y=-2182
XXB19A871F836 13 12 _GENERATED_158 _GENERATED_157 64 72 sram_filler $T=1152 -2182 0 0 $X=1156 $Y=-2182
XXB19A871F837 13 12 12 _GENERATED_159 64 72 sram_filler $T=816 -2182 0 0 $X=820 $Y=-2182
XXB19A871F838 13 12 _GENERATED_160 13 64 72 sram_filler $T=648 -2182 0 0 $X=652 $Y=-2182
XXB19A871F839 13 6 6 _GENERATED_161 64 71 sram_filler $T=1100 -2056 0 180 $X=652 $Y=-2646
XXB19A871F840 13 6 _GENERATED_162 13 64 71 sram_filler $T=1268 -2056 0 180 $X=820 $Y=-2646
XXB19A871F841 13 6 _GENERATED_164 _GENERATED_163 64 71 sram_filler $T=1604 -2056 0 180 $X=1156 $Y=-2646
XXB19A871F842 13 6 _GENERATED_166 _GENERATED_165 64 71 sram_filler $T=1940 -2056 0 180 $X=1492 $Y=-2646
XXB19A871F843 5 6 _GENERATED_168 _GENERATED_167 61 71 sram_filler $T=648 -3106 0 0 $X=652 $Y=-3106
XXB19A871F844 5 6 _GENERATED_170 _GENERATED_169 61 71 sram_filler $T=984 -3106 0 0 $X=988 $Y=-3106
XXB19A871F845 5 6 _GENERATED_171 5 61 71 sram_filler $T=1320 -3106 0 0 $X=1324 $Y=-3106
XXB19A871F846 5 6 6 _GENERATED_172 61 71 sram_filler $T=1488 -3106 0 0 $X=1492 $Y=-3106
XXB19A871F847 5 7 _GENERATED_174 _GENERATED_173 61 70 sram_filler $T=1940 -2980 0 180 $X=1492 $Y=-3570
XXB19A871F848 5 7 _GENERATED_176 _GENERATED_175 61 70 sram_filler $T=1604 -2980 0 180 $X=1156 $Y=-3570
XXB19A871F849 5 7 _GENERATED_177 5 61 70 sram_filler $T=1268 -2980 0 180 $X=820 $Y=-3570
XXB19A871F850 5 7 7 _GENERATED_178 61 70 sram_filler $T=1100 -2980 0 180 $X=652 $Y=-3570
XXB19A871F851 8 7 7 _GENERATED_179 62 70 sram_filler $T=1488 -4030 0 0 $X=1492 $Y=-4030
XXB19A871F852 8 7 _GENERATED_180 8 62 70 sram_filler $T=1320 -4030 0 0 $X=1324 $Y=-4030
XXB19A871F853 8 7 _GENERATED_182 _GENERATED_181 62 70 sram_filler $T=984 -4030 0 0 $X=988 $Y=-4030
XXB19A871F854 8 7 _GENERATED_184 _GENERATED_183 62 70 sram_filler $T=648 -4030 0 0 $X=652 $Y=-4030
XXB19A871F855 8 2 2 _GENERATED_185 62 69 sram_filler $T=1100 -3904 0 180 $X=652 $Y=-4494
XXB19A871F856 8 2 _GENERATED_186 8 62 69 sram_filler $T=1268 -3904 0 180 $X=820 $Y=-4494
XXB19A871F857 8 2 _GENERATED_188 _GENERATED_187 62 69 sram_filler $T=1604 -3904 0 180 $X=1156 $Y=-4494
XXB19A871F858 8 2 _GENERATED_190 _GENERATED_189 62 69 sram_filler $T=1940 -3904 0 180 $X=1492 $Y=-4494
XXB19A871F859 13 6 _GENERATED_192 _GENERATED_191 64 71 sram_filler $T=3168 -2056 1 0 $X=3172 $Y=-2646
XXB19A871F860 13 6 _GENERATED_194 _GENERATED_193 64 71 sram_filler $T=3840 -2056 1 0 $X=3844 $Y=-2646
XXB19A871F861 13 6 _GENERATED_196 _GENERATED_195 64 71 sram_filler $T=3504 -2056 1 0 $X=3508 $Y=-2646
XXB19A871F862 5 7 _GENERATED_198 _GENERATED_197 61 70 sram_filler $T=3840 -2980 1 0 $X=3844 $Y=-3570
XXB19A871F863 5 7 _GENERATED_200 _GENERATED_199 61 70 sram_filler $T=3168 -2980 1 0 $X=3172 $Y=-3570
XXB19A871F864 5 7 _GENERATED_202 _GENERATED_201 61 70 sram_filler $T=3504 -2980 1 0 $X=3508 $Y=-3570
XXB19A871F865 8 2 _GENERATED_204 _GENERATED_203 62 69 sram_filler $T=3168 -3904 1 0 $X=3172 $Y=-4494
XXB19A871F866 8 2 _GENERATED_206 _GENERATED_205 62 69 sram_filler $T=3840 -3904 1 0 $X=3844 $Y=-4494
XXB19A871F867 8 2 _GENERATED_208 _GENERATED_207 62 69 sram_filler $T=3504 -3904 1 0 $X=3508 $Y=-4494
XXB19A871F868 3 2 _GENERATED_210 _GENERATED_209 60 68 sram_filler $T=3840 -4828 1 0 $X=3844 $Y=-5418
XXB19A871F869 3 2 _GENERATED_212 _GENERATED_211 60 68 sram_filler $T=3168 -4828 1 0 $X=3172 $Y=-5418
XXB19A871F870 3 2 _GENERATED_214 _GENERATED_213 60 68 sram_filler $T=3504 -4828 1 0 $X=3508 $Y=-5418
XXB19A871F871 10 12 _GENERATED_216 _GENERATED_215 63 72 sram_filler $T=3504 -1132 1 0 $X=3508 $Y=-1722
XXB19A871F872 10 12 _GENERATED_218 _GENERATED_217 63 72 sram_filler $T=3168 -1132 1 0 $X=3172 $Y=-1722
XXB19A871F873 10 12 _GENERATED_220 _GENERATED_219 63 72 sram_filler $T=3840 -1132 1 0 $X=3844 $Y=-1722
XXB19A871F874 11 9 _GENERATED_222 _GENERATED_221 67 74 sram_filler $T=3504 -208 1 0 $X=3508 $Y=-798
XXB19A871F875 11 9 _GENERATED_224 _GENERATED_223 67 74 sram_filler $T=3840 -208 1 0 $X=3844 $Y=-798
XXB19A871F876 11 9 _GENERATED_226 _GENERATED_225 67 74 sram_filler $T=3168 -208 1 0 $X=3172 $Y=-798
XXB19A871F877 16 17 _GENERATED_228 _GENERATED_227 66 73 sram_filler $T=3168 716 1 0 $X=3172 $Y=126
XXB19A871F878 16 17 _GENERATED_230 _GENERATED_229 66 73 sram_filler $T=3840 716 1 0 $X=3844 $Y=126
XXB19A871F879 15 14 _GENERATED_232 _GENERATED_231 65 75 sram_filler $T=3840 1640 1 0 $X=3844 $Y=1050
XXB19A871F880 15 14 _GENERATED_234 _GENERATED_233 65 75 sram_filler $T=3168 1640 1 0 $X=3172 $Y=1050
XXB19A871F881 15 14 _GENERATED_236 _GENERATED_235 65 75 sram_filler $T=3504 1640 1 0 $X=3508 $Y=1050
XXB19A871F882 16 17 _GENERATED_238 _GENERATED_237 66 73 sram_filler $T=3504 716 1 0 $X=3508 $Y=126
XXB19A871F883 3 2 _GENERATED_240 _GENERATED_239 60 68 sram_filler $T=1488 -4828 1 0 $X=1492 $Y=-5418
XXB19A871F884 3 2 _GENERATED_242 _GENERATED_241 60 69 sram_filler $T=1488 -4954 0 0 $X=1492 $Y=-4954
.ends static_row_decoder_3by8
.subckt WLRef_PC 2 3 4 5 6 7 8 9 10 12 15
+	19 22 24 26 27 29 33 34 36 37 38
+	42 49 50 51 58 59 60 61 62 63 64
+	71
*.floating_nets 70
MM1 8 35 40 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5770 $Y=1241  $PIN_XY=5800,1136,5770,1241,5740,1136 $DEVICE_ID=1001
MM2 34 41 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5602 $Y=1661  $PIN_XY=5632,1766,5602,1661,5572,1766 $DEVICE_ID=1001
MM3 35 39 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5602 $Y=737  $PIN_XY=5632,842,5602,737,5572,842 $DEVICE_ID=1001
MM4 8 40 32 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5266 $Y=1241  $PIN_XY=5296,1136,5266,1241,5236,1136 $DEVICE_ID=1001
MM5 41 32 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5098 $Y=1661  $PIN_XY=5128,1766,5098,1661,5068,1766 $DEVICE_ID=1001
MM6 39 30 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5098 $Y=737  $PIN_XY=5128,842,5098,737,5068,842 $DEVICE_ID=1001
MM7 8 31 44 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4762 $Y=1241  $PIN_XY=4792,1136,4762,1241,4732,1136 $DEVICE_ID=1001
MM8 31 45 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4594 $Y=1682  $PIN_XY=4624,1766,4594,1682,4564,1766 $DEVICE_ID=1001
MM9 30 43 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4594 $Y=737  $PIN_XY=4624,842,4594,737,4564,842 $DEVICE_ID=1001
MM10 2 23 38 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4426 $Y=2165  $PIN_XY=4456,2060,4426,2165,4396,2060 $DEVICE_ID=1001
MM11 38 23 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4258 $Y=2165  $PIN_XY=4288,2060,4258,2165,4228,2060 $DEVICE_ID=1001
MM12 8 44 28 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4258 $Y=1241  $PIN_XY=4288,1136,4258,1241,4228,1136 $DEVICE_ID=1001
MM13 45 22 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4090 $Y=1661  $PIN_XY=4120,1766,4090,1661,4060,1766 $DEVICE_ID=1001
MM14 43 28 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4090 $Y=737  $PIN_XY=4120,842,4090,737,4060,842 $DEVICE_ID=1001
MM15 2 12 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3754 $Y=2144  $PIN_XY=3784,2060,3754,2144,3724,2060 $DEVICE_ID=1001
MM16 2 24 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3754 $Y=1703  $PIN_XY=3784,1766,3754,1703,3724,1766 $DEVICE_ID=1001
MM17 23 25 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3586 $Y=2165  $PIN_XY=3616,2060,3586,2165,3556,2060 $DEVICE_ID=1001
MM18 2 21 48 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3250 $Y=1661  $PIN_XY=3280,1766,3250,1661,3220,1766 $DEVICE_ID=1001
MM19 8 20 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3250 $Y=737  $PIN_XY=3280,842,3250,737,3220,842 $DEVICE_ID=1001
MM20 21 67 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3082 $Y=2144  $PIN_XY=3112,2060,3082,2144,3052,2060 $DEVICE_ID=1001
MM21 20 54 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3082 $Y=1241  $PIN_XY=3112,1136,3082,1241,3052,1136 $DEVICE_ID=1001
MM22 2 48 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2746 $Y=1661  $PIN_XY=2776,1766,2746,1661,2716,1766 $DEVICE_ID=1001
MM23 8 55 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2746 $Y=737  $PIN_XY=2776,842,2746,737,2716,842 $DEVICE_ID=1001
MM24 67 17 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2578 $Y=2144  $PIN_XY=2608,2060,2578,2144,2548,2060 $DEVICE_ID=1001
MM25 54 16 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2578 $Y=1241  $PIN_XY=2608,1136,2578,1241,2548,1136 $DEVICE_ID=1001
MM26 2 19 47 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2242 $Y=1661  $PIN_XY=2272,1766,2242,1661,2212,1766 $DEVICE_ID=1001
MM27 8 18 56 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2242 $Y=737  $PIN_XY=2272,842,2242,737,2212,842 $DEVICE_ID=1001
MM28 17 68 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2074 $Y=2144  $PIN_XY=2104,2060,2074,2144,2044,2060 $DEVICE_ID=1001
MM29 16 53 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2074 $Y=1241  $PIN_XY=2104,1136,2074,1241,2044,1136 $DEVICE_ID=1001
MM30 2 47 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1738 $Y=1661  $PIN_XY=1768,1766,1738,1661,1708,1766 $DEVICE_ID=1001
MM31 8 56 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1738 $Y=737  $PIN_XY=1768,842,1738,737,1708,842 $DEVICE_ID=1001
MM32 68 12 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1570 $Y=2144  $PIN_XY=1600,2060,1570,2144,1540,2060 $DEVICE_ID=1001
MM33 53 11 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1570 $Y=1241  $PIN_XY=1600,1136,1570,1241,1540,1136 $DEVICE_ID=1001
MM34 2 14 46 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1234 $Y=1661  $PIN_XY=1264,1766,1234,1661,1204,1766 $DEVICE_ID=1001
MM35 8 13 57 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1234 $Y=737  $PIN_XY=1264,842,1234,737,1204,842 $DEVICE_ID=1001
MM36 12 69 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1066 $Y=2144  $PIN_XY=1096,2060,1066,2144,1036,2060 $DEVICE_ID=1001
MM37 11 52 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1066 $Y=1241  $PIN_XY=1096,1136,1066,1241,1036,1136 $DEVICE_ID=1001
MM38 2 46 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=730 $Y=1661  $PIN_XY=760,1766,730,1661,700,1766 $DEVICE_ID=1001
MM39 8 57 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=730 $Y=737  $PIN_XY=760,842,730,737,700,842 $DEVICE_ID=1001
MM40 69 24 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=562 $Y=2144  $PIN_XY=592,2060,562,2144,532,2060 $DEVICE_ID=1001
MM41 52 25 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=562 $Y=1241  $PIN_XY=592,1136,562,1241,532,1136 $DEVICE_ID=1001
MM42 3 41 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5770 $Y=1581  $PIN_XY=5800,1596,5770,1581,5740,1596 $DEVICE_ID=1003
MM43 3 35 40 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5770 $Y=1241  $PIN_XY=5800,1306,5770,1241,5740,1306 $DEVICE_ID=1003
MM44 5 39 35 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5770 $Y=678  $PIN_XY=5800,672,5770,678,5740,672 $DEVICE_ID=1003
MM45 34 41 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5602 $Y=1661  $PIN_XY=5632,1596,5602,1661,5572,1596 $DEVICE_ID=1003
MM46 40 35 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5602 $Y=1321  $PIN_XY=5632,1306,5602,1321,5572,1306 $DEVICE_ID=1003
MM47 35 39 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5602 $Y=737  $PIN_XY=5632,672,5602,737,5572,672 $DEVICE_ID=1003
MM48 33 22 65 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5602 $Y=317  $PIN_XY=5632,382,5602,317,5572,382 $DEVICE_ID=1003
MM49 65 34 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5434 $Y=296  $PIN_XY=5464,382,5434,296,5404,382 $DEVICE_ID=1003
MM50 3 32 41 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5266 $Y=1581  $PIN_XY=5296,1596,5266,1581,5236,1596 $DEVICE_ID=1003
MM51 3 40 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5266 $Y=1241  $PIN_XY=5296,1306,5266,1241,5236,1306 $DEVICE_ID=1003
MM52 5 30 39 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5266 $Y=678  $PIN_XY=5296,672,5266,678,5236,672 $DEVICE_ID=1003
MM53 41 32 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5098 $Y=1661  $PIN_XY=5128,1596,5098,1661,5068,1596 $DEVICE_ID=1003
MM54 32 40 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5098 $Y=1321  $PIN_XY=5128,1306,5098,1321,5068,1306 $DEVICE_ID=1003
MM55 39 30 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5098 $Y=737  $PIN_XY=5128,672,5098,737,5068,672 $DEVICE_ID=1003
MM56 5 33 37 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5098 $Y=397  $PIN_XY=5128,382,5098,397,5068,382 $DEVICE_ID=1003
MM57 37 33 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4930 $Y=376  $PIN_XY=4960,382,4930,376,4900,382 $DEVICE_ID=1003
MM58 6 27 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=2585  $PIN_XY=4792,2520,4762,2585,4732,2520 $DEVICE_ID=1003
MM59 6 23 38 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=2245  $PIN_XY=4792,2230,4762,2245,4732,2230 $DEVICE_ID=1003
MM60 3 45 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=1581  $PIN_XY=4792,1596,4762,1581,4732,1596 $DEVICE_ID=1003
MM61 3 31 44 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=1241  $PIN_XY=4792,1306,4762,1241,4732,1306 $DEVICE_ID=1003
MM62 5 43 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4762 $Y=657  $PIN_XY=4792,672,4762,657,4732,672 $DEVICE_ID=1003
MM63 5 33 37 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4762 $Y=317  $PIN_XY=4792,382,4762,317,4732,382 $DEVICE_ID=1003
MM64 36 27 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4594 $Y=2585  $PIN_XY=4624,2520,4594,2585,4564,2520 $DEVICE_ID=1003
MM65 38 23 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4594 $Y=2245  $PIN_XY=4624,2230,4594,2245,4564,2230 $DEVICE_ID=1003
MM66 31 45 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4594 $Y=1682  $PIN_XY=4624,1596,4594,1682,4564,1596 $DEVICE_ID=1003
MM67 44 31 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4594 $Y=1321  $PIN_XY=4624,1306,4594,1321,4564,1306 $DEVICE_ID=1003
MM68 30 43 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4594 $Y=737  $PIN_XY=4624,672,4594,737,4564,672 $DEVICE_ID=1003
MM69 37 33 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4594 $Y=317  $PIN_XY=4624,382,4594,317,4564,382 $DEVICE_ID=1003
MM70 6 27 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4426 $Y=2505  $PIN_XY=4456,2520,4426,2505,4396,2520 $DEVICE_ID=1003
MM71 6 23 38 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4426 $Y=2165  $PIN_XY=4456,2230,4426,2165,4396,2230 $DEVICE_ID=1003
MM72 36 27 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4258 $Y=2505  $PIN_XY=4288,2520,4258,2505,4228,2520 $DEVICE_ID=1003
MM73 38 23 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4258 $Y=2165  $PIN_XY=4288,2230,4258,2165,4228,2230 $DEVICE_ID=1003
MM74 3 22 45 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4258 $Y=1581  $PIN_XY=4288,1596,4258,1581,4228,1596 $DEVICE_ID=1003
MM75 3 44 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4258 $Y=1241  $PIN_XY=4288,1306,4258,1241,4228,1306 $DEVICE_ID=1003
MM76 5 28 43 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4258 $Y=657  $PIN_XY=4288,672,4258,657,4228,672 $DEVICE_ID=1003
MM77 5 42 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4258 $Y=397  $PIN_XY=4288,382,4258,397,4228,382 $DEVICE_ID=1003
MM78 45 22 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4090 $Y=1661  $PIN_XY=4120,1596,4090,1661,4060,1596 $DEVICE_ID=1003
MM79 28 44 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4090 $Y=1321  $PIN_XY=4120,1306,4090,1321,4060,1306 $DEVICE_ID=1003
MM80 43 28 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4090 $Y=737  $PIN_XY=4120,672,4090,737,4060,672 $DEVICE_ID=1003
MM81 29 42 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4090 $Y=317  $PIN_XY=4120,382,4090,317,4060,382 $DEVICE_ID=1003
MM82 6 19 27 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3754 $Y=2585  $PIN_XY=3784,2520,3754,2585,3724,2520 $DEVICE_ID=1003
MM83 23 12 66 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3754 $Y=2144  $PIN_XY=3784,2230,3754,2144,3724,2230 $DEVICE_ID=1003
MM84 3 24 22 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3754 $Y=1703  $PIN_XY=3784,1596,3754,1703,3724,1596 $DEVICE_ID=1003
MM85 5 26 42 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3754 $Y=376  $PIN_XY=3784,382,3754,376,3724,382 $DEVICE_ID=1003
MM86 27 12 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3586 $Y=2585  $PIN_XY=3616,2520,3586,2585,3556,2520 $DEVICE_ID=1003
MM87 66 25 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3586 $Y=2165  $PIN_XY=3616,2230,3586,2165,3556,2230 $DEVICE_ID=1003
MM88 22 24 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3586 $Y=1602  $PIN_XY=3616,1596,3586,1602,3556,1596 $DEVICE_ID=1003
MM89 42 26 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3586 $Y=296  $PIN_XY=3616,382,3586,296,3556,382 $DEVICE_ID=1003
MM90 6 67 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3250 $Y=2224  $PIN_XY=3280,2230,3250,2224,3220,2230 $DEVICE_ID=1003
MM91 3 21 48 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3250 $Y=1661  $PIN_XY=3280,1596,3250,1661,3220,1596 $DEVICE_ID=1003
MM92 3 54 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3250 $Y=1321  $PIN_XY=3280,1306,3250,1321,3220,1306 $DEVICE_ID=1003
MM93 5 20 55 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3250 $Y=737  $PIN_XY=3280,672,3250,737,3220,672 $DEVICE_ID=1003
MM94 5 51 26 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3250 $Y=397  $PIN_XY=3280,382,3250,397,3220,382 $DEVICE_ID=1003
MM95 21 67 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3082 $Y=2144  $PIN_XY=3112,2230,3082,2144,3052,2230 $DEVICE_ID=1003
MM96 48 21 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3082 $Y=1581  $PIN_XY=3112,1596,3082,1581,3052,1596 $DEVICE_ID=1003
MM97 20 54 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3082 $Y=1241  $PIN_XY=3112,1306,3082,1241,3052,1306 $DEVICE_ID=1003
MM98 55 20 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3082 $Y=657  $PIN_XY=3112,672,3082,657,3052,672 $DEVICE_ID=1003
MM99 26 51 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3082 $Y=317  $PIN_XY=3112,382,3082,317,3052,382 $DEVICE_ID=1003
MM100 6 17 67 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2746 $Y=2224  $PIN_XY=2776,2230,2746,2224,2716,2230 $DEVICE_ID=1003
MM101 3 48 19 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2746 $Y=1661  $PIN_XY=2776,1596,2746,1661,2716,1596 $DEVICE_ID=1003
MM102 3 16 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2746 $Y=1321  $PIN_XY=2776,1306,2746,1321,2716,1306 $DEVICE_ID=1003
MM103 5 55 18 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2746 $Y=737  $PIN_XY=2776,672,2746,737,2716,672 $DEVICE_ID=1003
MM104 5 15 51 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2746 $Y=397  $PIN_XY=2776,382,2746,397,2716,382 $DEVICE_ID=1003
MM105 67 17 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2578 $Y=2144  $PIN_XY=2608,2230,2578,2144,2548,2230 $DEVICE_ID=1003
MM106 19 48 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2578 $Y=1581  $PIN_XY=2608,1596,2578,1581,2548,1596 $DEVICE_ID=1003
MM107 54 16 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2578 $Y=1241  $PIN_XY=2608,1306,2578,1241,2548,1306 $DEVICE_ID=1003
MM108 18 55 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2578 $Y=657  $PIN_XY=2608,672,2578,657,2548,672 $DEVICE_ID=1003
MM109 51 15 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2578 $Y=317  $PIN_XY=2608,382,2578,317,2548,382 $DEVICE_ID=1003
MM110 6 68 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2242 $Y=2224  $PIN_XY=2272,2230,2242,2224,2212,2230 $DEVICE_ID=1003
MM111 3 19 47 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2242 $Y=1661  $PIN_XY=2272,1596,2242,1661,2212,1596 $DEVICE_ID=1003
MM112 3 53 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2242 $Y=1321  $PIN_XY=2272,1306,2242,1321,2212,1306 $DEVICE_ID=1003
MM113 5 18 56 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2242 $Y=737  $PIN_XY=2272,672,2242,737,2212,672 $DEVICE_ID=1003
MM114 5 50 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2242 $Y=397  $PIN_XY=2272,382,2242,397,2212,382 $DEVICE_ID=1003
MM115 17 68 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2074 $Y=2144  $PIN_XY=2104,2230,2074,2144,2044,2230 $DEVICE_ID=1003
MM116 47 19 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2074 $Y=1581  $PIN_XY=2104,1596,2074,1581,2044,1596 $DEVICE_ID=1003
MM117 16 53 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2074 $Y=1241  $PIN_XY=2104,1306,2074,1241,2044,1306 $DEVICE_ID=1003
MM118 56 18 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2074 $Y=657  $PIN_XY=2104,672,2074,657,2044,672 $DEVICE_ID=1003
MM119 15 50 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2074 $Y=317  $PIN_XY=2104,382,2074,317,2044,382 $DEVICE_ID=1003
MM120 6 12 68 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1738 $Y=2224  $PIN_XY=1768,2230,1738,2224,1708,2230 $DEVICE_ID=1003
MM121 3 47 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1738 $Y=1661  $PIN_XY=1768,1596,1738,1661,1708,1596 $DEVICE_ID=1003
MM122 3 11 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1738 $Y=1321  $PIN_XY=1768,1306,1738,1321,1708,1306 $DEVICE_ID=1003
MM123 5 56 13 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1738 $Y=737  $PIN_XY=1768,672,1738,737,1708,672 $DEVICE_ID=1003
MM124 5 10 50 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1738 $Y=397  $PIN_XY=1768,382,1738,397,1708,382 $DEVICE_ID=1003
MM125 68 12 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1570 $Y=2144  $PIN_XY=1600,2230,1570,2144,1540,2230 $DEVICE_ID=1003
MM126 14 47 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1570 $Y=1581  $PIN_XY=1600,1596,1570,1581,1540,1596 $DEVICE_ID=1003
MM127 53 11 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1570 $Y=1241  $PIN_XY=1600,1306,1570,1241,1540,1306 $DEVICE_ID=1003
MM128 13 56 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1570 $Y=657  $PIN_XY=1600,672,1570,657,1540,672 $DEVICE_ID=1003
MM129 50 10 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1570 $Y=317  $PIN_XY=1600,382,1570,317,1540,382 $DEVICE_ID=1003
MM130 6 69 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1234 $Y=2224  $PIN_XY=1264,2230,1234,2224,1204,2230 $DEVICE_ID=1003
MM131 3 14 46 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1234 $Y=1661  $PIN_XY=1264,1596,1234,1661,1204,1596 $DEVICE_ID=1003
MM132 3 52 11 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1234 $Y=1321  $PIN_XY=1264,1306,1234,1321,1204,1306 $DEVICE_ID=1003
MM133 5 13 57 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1234 $Y=737  $PIN_XY=1264,672,1234,737,1204,672 $DEVICE_ID=1003
MM134 5 49 10 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1234 $Y=397  $PIN_XY=1264,382,1234,397,1204,382 $DEVICE_ID=1003
MM135 12 69 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1066 $Y=2144  $PIN_XY=1096,2230,1066,2144,1036,2230 $DEVICE_ID=1003
MM136 46 14 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1066 $Y=1581  $PIN_XY=1096,1596,1066,1581,1036,1596 $DEVICE_ID=1003
MM137 11 52 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1066 $Y=1241  $PIN_XY=1096,1306,1066,1241,1036,1306 $DEVICE_ID=1003
MM138 57 13 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1066 $Y=657  $PIN_XY=1096,672,1066,657,1036,672 $DEVICE_ID=1003
MM139 10 49 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1066 $Y=317  $PIN_XY=1096,382,1066,317,1036,382 $DEVICE_ID=1003
MM140 6 24 69 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=730 $Y=2224  $PIN_XY=760,2230,730,2224,700,2230 $DEVICE_ID=1003
MM141 3 46 25 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=730 $Y=1661  $PIN_XY=760,1596,730,1661,700,1596 $DEVICE_ID=1003
MM142 3 25 52 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=730 $Y=1321  $PIN_XY=760,1306,730,1321,700,1306 $DEVICE_ID=1003
MM143 5 57 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=730 $Y=737  $PIN_XY=760,672,730,737,700,672 $DEVICE_ID=1003
MM144 5 9 49 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=730 $Y=397  $PIN_XY=760,382,730,397,700,382 $DEVICE_ID=1003
MM145 69 24 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=562 $Y=2144  $PIN_XY=592,2230,562,2144,532,2230 $DEVICE_ID=1003
MM146 25 46 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=562 $Y=1581  $PIN_XY=592,1596,562,1581,532,1596 $DEVICE_ID=1003
MM147 52 25 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=562 $Y=1241  $PIN_XY=592,1306,562,1241,532,1306 $DEVICE_ID=1003
MM148 9 57 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=562 $Y=657  $PIN_XY=592,672,562,657,532,672 $DEVICE_ID=1003
MM149 49 9 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=562 $Y=317  $PIN_XY=592,382,562,317,532,382 $DEVICE_ID=1003
XXB19A871F885 2 3 22 24 59 62 inv $T=3976 1976 0 180 $X=3364 $Y=1386
XXB19A871F886 4 5 33 22 34 65 61 63 nor $T=4584 0 0 0 $X=5212 $Y=2
XXB19A871F887 2 6 23 12 25 66 59 64 nor $T=2736 1848 0 0 $X=3364 $Y=1850
XXB19A871F888 7 6 27 12 19 71 58 64 nand $T=2946 3128 1 0 $X=3364 $Y=2310
XXB19A871F889 7 6 36 27 58 64 invx4 $T=5008 2900 0 180 $X=4035 $Y=2310
XXB19A871F890 4 5 37 33 61 63 invx4 $T=4348 2 0 0 $X=4372 $Y=2
XXB19A871F891 2 6 38 23 59 64 invx4 $T=4012 1850 0 0 $X=4036 $Y=1850
XXB19A871F892 8 5 39 35 30 60 63 buffer $T=4796 1054 1 0 $X=4876 $Y=462
XXB19A871F893 8 3 40 32 35 60 62 buffer $T=6072 924 1 180 $X=4876 $Y=926
XXB19A871F894 2 3 41 34 32 59 62 buffer $T=4796 1978 1 0 $X=4876 $Y=1386
XXB19A871F895 4 5 42 29 26 61 63 buffer $T=3284 0 0 0 $X=3364 $Y=2
XXB19A871F896 8 5 43 30 28 60 63 buffer $T=3788 1054 1 0 $X=3868 $Y=462
XXB19A871F897 8 3 44 28 31 60 62 buffer $T=5064 924 1 180 $X=3868 $Y=926
XXB19A871F898 2 3 45 31 22 59 62 buffer $T=3788 1978 1 0 $X=3868 $Y=1386
XXB19A871F899 2 3 46 25 14 59 62 buffer $T=1536 1978 0 180 $X=340 $Y=1386
XXB19A871F900 2 3 47 14 19 59 62 buffer $T=2544 1978 0 180 $X=1348 $Y=1386
XXB19A871F901 2 3 48 19 21 59 62 buffer $T=3552 1978 0 180 $X=2356 $Y=1386
XXB19A871F902 2 6 67 21 17 59 64 buffer $T=2276 1848 0 0 $X=2356 $Y=1850
XXB19A871F903 2 6 68 17 12 59 64 buffer $T=1268 1848 0 0 $X=1348 $Y=1850
XXB19A871F904 2 6 69 12 24 59 64 buffer $T=260 1848 0 0 $X=340 $Y=1850
XXB19A871F905 4 5 49 10 9 61 63 buffer $T=260 0 0 0 $X=340 $Y=2
XXB19A871F906 4 5 50 15 10 61 63 buffer $T=1268 0 0 0 $X=1348 $Y=2
XXB19A871F907 4 5 51 26 15 61 63 buffer $T=2276 0 0 0 $X=2356 $Y=2
XXB19A871F908 8 3 52 11 25 60 62 buffer $T=260 924 0 0 $X=340 $Y=926
XXB19A871F909 8 3 53 16 11 60 62 buffer $T=1268 924 0 0 $X=1348 $Y=926
XXB19A871F910 8 3 54 20 16 60 62 buffer $T=2276 924 0 0 $X=2356 $Y=926
XXB19A871F911 8 5 55 18 20 60 63 buffer $T=3552 1054 0 180 $X=2356 $Y=462
XXB19A871F912 8 5 56 13 18 60 63 buffer $T=2544 1054 0 180 $X=1348 $Y=462
XXB19A871F913 8 5 57 9 13 60 63 buffer $T=1536 1054 0 180 $X=340 $Y=462
XXB19A871F914 7 6 _GENERATED_73 _GENERATED_72 58 64 sram_filler $T=788 2900 0 180 $X=340 $Y=2310
XXB19A871F915 7 6 _GENERATED_75 _GENERATED_74 58 64 sram_filler $T=1124 2900 0 180 $X=676 $Y=2310
XXB19A871F916 7 6 _GENERATED_77 _GENERATED_76 58 64 sram_filler $T=1460 2900 0 180 $X=1012 $Y=2310
XXB19A871F917 7 6 _GENERATED_79 _GENERATED_78 58 64 sram_filler $T=1796 2900 0 180 $X=1348 $Y=2310
XXB19A871F918 7 6 _GENERATED_81 _GENERATED_80 58 64 sram_filler $T=2132 2900 0 180 $X=1684 $Y=2310
XXB19A871F919 7 6 _GENERATED_83 _GENERATED_82 58 64 sram_filler $T=2468 2900 0 180 $X=2020 $Y=2310
XXB19A871F920 7 6 _GENERATED_85 _GENERATED_84 58 64 sram_filler $T=2804 2900 0 180 $X=2356 $Y=2310
XXB19A871F921 7 6 _GENERATED_87 _GENERATED_86 58 64 sram_filler $T=3140 2900 0 180 $X=2692 $Y=2310
XXB19A871F922 7 6 _GENERATED_89 _GENERATED_88 58 64 sram_filler $T=3476 2900 0 180 $X=3028 $Y=2310
XXB19A871F923 7 6 _GENERATED_91 _GENERATED_90 58 64 sram_filler $T=5996 2900 0 180 $X=5548 $Y=2310
XXB19A871F924 7 6 _GENERATED_93 _GENERATED_92 58 64 sram_filler $T=5660 2900 0 180 $X=5212 $Y=2310
XXB19A871F925 7 6 _GENERATED_95 _GENERATED_94 58 64 sram_filler $T=5324 2900 0 180 $X=4875 $Y=2310
XXB19A871F926 2 6 _GENERATED_97 _GENERATED_96 59 64 sram_filler $T=5544 1850 0 0 $X=5548 $Y=1850
XXB19A871F927 2 6 _GENERATED_99 _GENERATED_98 59 64 sram_filler $T=5208 1850 0 0 $X=5212 $Y=1850
XXB19A871F928 2 6 _GENERATED_101 _GENERATED_100 59 64 sram_filler $T=4872 1850 0 0 $X=4875 $Y=1850
XXB19A871F929 8 5 5 _GENERATED_102 60 63 sram_filler $T=3812 1052 0 180 $X=3364 $Y=462
XXB19A871F930 8 5 _GENERATED_103 8 60 63 sram_filler $T=3980 1052 0 180 $X=3532 $Y=462
XXB19A871F931 8 3 3 _GENERATED_104 60 62 sram_filler $T=3528 926 0 0 $X=3532 $Y=926
XXB19A871F932 8 3 _GENERATED_105 8 60 62 sram_filler $T=3360 926 0 0 $X=3364 $Y=926
.ends WLRef_PC
.subckt agen_unit 2 3 4 5 6 7 8 9 10 14 15
+	18 19 20 23 26 27 28 29 30 31 32
+	33 35 37 38 39 40 41 42 43 44 45
+	46 47 59 60 61
MM1 8 23 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=1895  $PIN_XY=3782,1832,3752,1895,3722,1832 $DEVICE_ID=1001
MM2 8 25 26 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=1454  $PIN_XY=3782,1538,3752,1454,3722,1538 $DEVICE_ID=1001
MM3 10 21 32 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=992  $PIN_XY=3782,908,3752,992,3722,908 $DEVICE_ID=1001
MM4 10 36 31 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=530  $PIN_XY=3782,614,3752,530,3722,614 $DEVICE_ID=1001
MM5 3 24 30 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=68  $PIN_XY=3782,-16,3752,68,3722,-16 $DEVICE_ID=1001
MM6 3 22 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=-394  $PIN_XY=3782,-310,3752,-394,3722,-310 $DEVICE_ID=1001
MM7 5 34 28 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=-856  $PIN_XY=3782,-940,3752,-856,3722,-940 $DEVICE_ID=1001
MM8 5 35 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=-1297  $PIN_XY=3782,-1234,3752,-1297,3722,-1234 $DEVICE_ID=1001
MM9 33 23 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=1895  $PIN_XY=3614,1832,3584,1895,3554,1832 $DEVICE_ID=1001
MM10 26 25 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=1454  $PIN_XY=3614,1538,3584,1454,3554,1538 $DEVICE_ID=1001
MM11 32 21 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=992  $PIN_XY=3614,908,3584,992,3554,908 $DEVICE_ID=1001
MM12 31 36 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=530  $PIN_XY=3614,614,3584,530,3554,614 $DEVICE_ID=1001
MM13 30 24 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=68  $PIN_XY=3614,-16,3584,68,3554,-16 $DEVICE_ID=1001
MM14 29 22 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-394  $PIN_XY=3614,-310,3584,-394,3554,-310 $DEVICE_ID=1001
MM15 28 34 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-856  $PIN_XY=3614,-940,3584,-856,3554,-940 $DEVICE_ID=1001
MM16 27 35 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-1297  $PIN_XY=3614,-1234,3584,-1297,3554,-1234 $DEVICE_ID=1001
MM17 10 12 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=971  $PIN_XY=3278,908,3248,971,3218,908 $DEVICE_ID=1001
MM18 10 17 36 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=551  $PIN_XY=3278,614,3248,551,3218,614 $DEVICE_ID=1001
MM19 5 11 34 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=-877  $PIN_XY=3278,-940,3248,-877,3218,-940 $DEVICE_ID=1001
MM20 5 15 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=-1297  $PIN_XY=3278,-1234,3248,-1297,3218,-1234 $DEVICE_ID=1001
MM21 23 20 58 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=1895  $PIN_XY=3110,1832,3080,1895,3050,1832 $DEVICE_ID=1001
MM22 25 20 57 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=1454  $PIN_XY=3110,1538,3080,1454,3050,1538 $DEVICE_ID=1001
MM23 21 20 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=992  $PIN_XY=3110,908,3080,992,3050,908 $DEVICE_ID=1001
MM24 36 20 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=530  $PIN_XY=3110,614,3080,530,3050,614 $DEVICE_ID=1001
MM25 24 20 56 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=68  $PIN_XY=3110,-16,3080,68,3050,-16 $DEVICE_ID=1001
MM26 22 20 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=-394  $PIN_XY=3110,-310,3080,-394,3050,-310 $DEVICE_ID=1001
MM27 34 20 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=-856  $PIN_XY=3110,-940,3080,-856,3050,-940 $DEVICE_ID=1001
MM28 35 20 5 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=-1297  $PIN_XY=3110,-1234,3080,-1297,3050,-1234 $DEVICE_ID=1001
MM29 58 18 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=1895  $PIN_XY=2942,1832,2912,1895,2882,1832 $DEVICE_ID=1001
MM30 57 14 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=1475  $PIN_XY=2942,1538,2912,1475,2882,1538 $DEVICE_ID=1001
MM31 56 16 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=47  $PIN_XY=2942,-16,2912,47,2882,-16 $DEVICE_ID=1001
MM32 55 13 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=-373  $PIN_XY=2942,-310,2912,-373,2882,-310 $DEVICE_ID=1001
MM33 20 19 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2408 $Y=992  $PIN_XY=2438,908,2408,992,2378,908 $DEVICE_ID=1001
MM34 8 12 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2072 $Y=1454  $PIN_XY=2102,1538,2072,1454,2042,1538 $DEVICE_ID=1001
MM35 3 11 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2072 $Y=-394  $PIN_XY=2102,-310,2072,-394,2042,-310 $DEVICE_ID=1001
MM36 18 14 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1904 $Y=1916  $PIN_XY=1934,1832,1904,1916,1874,1832 $DEVICE_ID=1001
MM37 16 13 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1904 $Y=68  $PIN_XY=1934,-16,1904,68,1874,-16 $DEVICE_ID=1001
MM38 7 25 26 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=1353  $PIN_XY=4118,1368,4088,1353,4058,1368 $DEVICE_ID=1003
MM39 7 21 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=1093  $PIN_XY=4118,1078,4088,1093,4058,1078 $DEVICE_ID=1003
MM40 4 36 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=429  $PIN_XY=4118,444,4088,429,4058,444 $DEVICE_ID=1003
MM41 4 24 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=169  $PIN_XY=4118,154,4088,169,4058,154 $DEVICE_ID=1003
MM42 2 22 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=-495  $PIN_XY=4118,-480,4088,-495,4058,-480 $DEVICE_ID=1003
MM43 2 34 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=-755  $PIN_XY=4118,-770,4088,-755,4058,-770 $DEVICE_ID=1003
MM44 26 25 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=1353  $PIN_XY=3950,1368,3920,1353,3890,1368 $DEVICE_ID=1003
MM45 32 21 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=1093  $PIN_XY=3950,1078,3920,1093,3890,1078 $DEVICE_ID=1003
MM46 31 36 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=429  $PIN_XY=3950,444,3920,429,3890,444 $DEVICE_ID=1003
MM47 30 24 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=169  $PIN_XY=3950,154,3920,169,3890,154 $DEVICE_ID=1003
MM48 29 22 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=-495  $PIN_XY=3950,-480,3920,-495,3890,-480 $DEVICE_ID=1003
MM49 28 34 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=-755  $PIN_XY=3950,-770,3920,-755,3890,-770 $DEVICE_ID=1003
MM50 7 25 26 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=1454  $PIN_XY=3782,1368,3752,1454,3722,1368 $DEVICE_ID=1003
MM51 7 21 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=992  $PIN_XY=3782,1078,3752,992,3722,1078 $DEVICE_ID=1003
MM52 4 36 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=530  $PIN_XY=3782,444,3752,530,3722,444 $DEVICE_ID=1003
MM53 4 24 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=68  $PIN_XY=3782,154,3752,68,3722,154 $DEVICE_ID=1003
MM54 2 22 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=-394  $PIN_XY=3782,-480,3752,-394,3722,-480 $DEVICE_ID=1003
MM55 2 34 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=-856  $PIN_XY=3782,-770,3752,-856,3722,-770 $DEVICE_ID=1003
MM56 26 25 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=1454  $PIN_XY=3614,1368,3584,1454,3554,1368 $DEVICE_ID=1003
MM57 32 21 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=992  $PIN_XY=3614,1078,3584,992,3554,1078 $DEVICE_ID=1003
MM58 31 36 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=530  $PIN_XY=3614,444,3584,530,3554,444 $DEVICE_ID=1003
MM59 30 24 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=68  $PIN_XY=3614,154,3584,68,3554,154 $DEVICE_ID=1003
MM60 29 22 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-394  $PIN_XY=3614,-480,3584,-394,3554,-480 $DEVICE_ID=1003
MM61 28 34 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-856  $PIN_XY=3614,-770,3584,-856,3554,-770 $DEVICE_ID=1003
MM62 7 12 50 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=971  $PIN_XY=3278,1078,3248,971,3218,1078 $DEVICE_ID=1003
MM63 4 17 49 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=551  $PIN_XY=3278,444,3248,551,3218,444 $DEVICE_ID=1003
MM64 2 11 48 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=-877  $PIN_XY=3278,-770,3248,-877,3218,-770 $DEVICE_ID=1003
MM65 7 20 25 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=1454  $PIN_XY=3110,1368,3080,1454,3050,1368 $DEVICE_ID=1003
MM66 50 20 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=992  $PIN_XY=3110,1078,3080,992,3050,1078 $DEVICE_ID=1003
MM67 49 20 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=530  $PIN_XY=3110,444,3080,530,3050,444 $DEVICE_ID=1003
MM68 4 20 24 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=68  $PIN_XY=3110,154,3080,68,3050,154 $DEVICE_ID=1003
MM69 2 20 22 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=-394  $PIN_XY=3110,-480,3080,-394,3050,-480 $DEVICE_ID=1003
MM70 48 20 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=-856  $PIN_XY=3110,-770,3080,-856,3050,-770 $DEVICE_ID=1003
MM71 25 14 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=1475  $PIN_XY=2942,1368,2912,1475,2882,1368 $DEVICE_ID=1003
MM72 24 16 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=47  $PIN_XY=2942,154,2912,47,2882,154 $DEVICE_ID=1003
MM73 22 13 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=-373  $PIN_XY=2942,-480,2912,-373,2882,-480 $DEVICE_ID=1003
MM74 7 19 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2576 $Y=1072  $PIN_XY=2606,1078,2576,1072,2546,1078 $DEVICE_ID=1003
MM75 20 19 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2408 $Y=992  $PIN_XY=2438,1078,2408,992,2378,1078 $DEVICE_ID=1003
MM76 7 12 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2072 $Y=1454  $PIN_XY=2102,1368,2072,1454,2042,1368 $DEVICE_ID=1003
MM77 4 13 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2072 $Y=154  $PIN_XY=2102,154,2072,154,2042,154 $DEVICE_ID=1003
MM78 2 11 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2072 $Y=-394  $PIN_XY=2102,-480,2072,-394,2042,-480 $DEVICE_ID=1003
MM79 17 12 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1904 $Y=1374  $PIN_XY=1934,1368,1904,1374,1874,1368 $DEVICE_ID=1003
MM80 16 13 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1904 $Y=68  $PIN_XY=1934,154,1904,68,1874,154 $DEVICE_ID=1003
MM81 15 11 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1904 $Y=-474  $PIN_XY=1934,-480,1904,-474,1874,-480 $DEVICE_ID=1003
MM82 7 54 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1568 $Y=1374  $PIN_XY=1598,1368,1568,1374,1538,1368 $DEVICE_ID=1003
MM83 4 52 13 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1568 $Y=148  $PIN_XY=1598,154,1568,148,1538,154 $DEVICE_ID=1003
MM84 2 53 11 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1568 $Y=-474  $PIN_XY=1598,-480,1568,-474,1538,-480 $DEVICE_ID=1003
MM85 12 54 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1400 $Y=1475  $PIN_XY=1430,1368,1400,1475,1370,1368 $DEVICE_ID=1003
MM86 13 52 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1400 $Y=47  $PIN_XY=1430,154,1400,47,1370,154 $DEVICE_ID=1003
MM87 11 53 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1400 $Y=-373  $PIN_XY=1430,-480,1400,-373,1370,-480 $DEVICE_ID=1003
MM88 7 19 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=896 $Y=1475  $PIN_XY=926,1368,896,1475,866,1368 $DEVICE_ID=1003
MM89 4 51 52 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=896 $Y=47  $PIN_XY=926,154,896,47,866,154 $DEVICE_ID=1003
MM90 2 19 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=896 $Y=-373  $PIN_XY=926,-480,896,-373,866,-480 $DEVICE_ID=1003
MM91 54 38 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=728 $Y=1475  $PIN_XY=758,1368,728,1475,698,1368 $DEVICE_ID=1003
MM92 52 37 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=728 $Y=47  $PIN_XY=758,154,728,47,698,154 $DEVICE_ID=1003
MM93 53 37 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=728 $Y=-373  $PIN_XY=758,-480,728,-373,698,-480 $DEVICE_ID=1003
MM94 4 19 51 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=392 $Y=148  $PIN_XY=422,154,392,148,362,154 $DEVICE_ID=1003
MM95 51 19 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=224 $Y=68  $PIN_XY=254,154,224,68,194,154 $DEVICE_ID=1003
XXB19A871F933 3 2 15 11 41 43 inv $T=2294 -100 0 180 $X=1682 $Y=-690
XXB19A871F934 3 4 16 13 41 44 inv $T=1682 -226 0 0 $X=1682 $Y=-226
XXB19A871F935 10 7 20 19 40 46 inv $T=2186 698 0 0 $X=2186 $Y=698
XXB19A871F936 8 7 17 12 42 46 inv $T=2294 1748 0 180 $X=1682 $Y=1158
XXB19A871F937 8 9 18 14 42 47 inv $T=1682 1622 0 0 $X=1682 $Y=1622
XXB19A871F938 5 2 34 20 11 48 39 43 nor $T=4098 -1152 1 180 $X=2690 $Y=-1150
XXB19A871F939 5 6 35 20 15 59 39 45 nor $T=4098 -1022 0 180 $X=2690 $Y=-1613
XXB19A871F940 10 4 36 20 17 49 40 44 nor $T=4098 826 0 180 $X=2690 $Y=234
XXB19A871F941 10 7 21 20 12 50 40 46 nor $T=4098 696 1 180 $X=2690 $Y=698
XXB19A871F942 3 2 22 13 20 55 41 43 nand $T=2272 128 1 0 $X=2690 $Y=-690
XXB19A871F943 3 4 24 16 20 56 41 44 nand $T=2272 -454 0 0 $X=2690 $Y=-226
XXB19A871F944 8 7 25 14 20 57 42 46 nand $T=2272 1976 1 0 $X=2690 $Y=1158
XXB19A871F945 8 9 23 18 20 58 42 47 nand $T=2272 1394 0 0 $X=2690 $Y=1622
XXB19A871F946 3 2 4 19 51 37 53 52 11 13 41 
+	43 44 Demux $T=2 -688 0 0 $X=2 $Y=-690
XXB19A871F947 8 7 9 19 60 38 54 61 12 14 42 
+	46 47 Demux $T=2 1160 0 0 $X=2 $Y=1158
XXB19A871F948 3 4 30 24 41 44 invx4 $T=3338 -226 0 0 $X=3362 $Y=-226
XXB19A871F949 10 4 31 36 40 44 invx4 $T=3338 824 1 0 $X=3362 $Y=234
XXB19A871F950 5 6 27 35 39 45 invx4 $T=3338 -1024 1 0 $X=3362 $Y=-1613
XXB19A871F951 3 2 29 22 41 43 invx4 $T=3338 -100 1 0 $X=3362 $Y=-690
XXB19A871F952 5 2 28 34 39 43 invx4 $T=3338 -1150 0 0 $X=3362 $Y=-1150
XXB19A871F953 8 9 33 23 42 47 invx4 $T=3338 1622 0 0 $X=3362 $Y=1622
XXB19A871F954 8 7 26 25 42 46 invx4 $T=3338 1748 1 0 $X=3362 $Y=1158
XXB19A871F955 10 7 32 21 40 46 invx4 $T=3338 698 0 0 $X=3362 $Y=698
XXB19A871F956 5 6 _GENERATED_63 _GENERATED_62 39 45 sram_filler $T=-2 -1024 1 0 $X=2 $Y=-1613
XXB19A871F957 5 6 _GENERATED_64 5 39 45 sram_filler $T=334 -1024 1 0 $X=338 $Y=-1613
XXB19A871F958 5 6 6 _GENERATED_65 39 45 sram_filler $T=502 -1024 1 0 $X=506 $Y=-1613
XXB19A871F959 5 2 _GENERATED_66 5 39 43 sram_filler $T=-2 -1150 0 0 $X=2 $Y=-1150
XXB19A871F960 5 2 2 _GENERATED_67 39 43 sram_filler $T=166 -1150 0 0 $X=170 $Y=-1150
XXB19A871F961 5 2 _GENERATED_69 _GENERATED_68 39 43 sram_filler $T=502 -1150 0 0 $X=506 $Y=-1150
XXB19A871F962 5 6 6 _GENERATED_70 39 45 sram_filler $T=1342 -1024 1 0 $X=1346 $Y=-1613
XXB19A871F963 5 6 _GENERATED_71 5 39 45 sram_filler $T=1174 -1024 1 0 $X=1178 $Y=-1613
XXB19A871F964 5 6 _GENERATED_73 _GENERATED_72 39 45 sram_filler $T=838 -1024 1 0 $X=842 $Y=-1613
XXB19A871F965 5 2 2 _GENERATED_74 39 43 sram_filler $T=1342 -1150 0 0 $X=1346 $Y=-1150
XXB19A871F966 5 2 _GENERATED_75 5 39 43 sram_filler $T=1174 -1150 0 0 $X=1178 $Y=-1150
XXB19A871F967 5 2 _GENERATED_77 _GENERATED_76 39 43 sram_filler $T=838 -1150 0 0 $X=842 $Y=-1150
XXB19A871F968 5 2 _GENERATED_79 _GENERATED_78 39 43 sram_filler $T=1678 -1150 0 0 $X=1682 $Y=-1150
XXB19A871F969 5 6 _GENERATED_81 _GENERATED_80 39 45 sram_filler $T=2130 -1024 0 180 $X=1682 $Y=-1613
XXB19A871F970 10 7 7 _GENERATED_82 40 46 sram_filler $T=1846 698 0 0 $X=1850 $Y=698
XXB19A871F971 10 4 _GENERATED_83 10 40 44 sram_filler $T=2298 824 0 180 $X=1850 $Y=234
XXB19A871F972 5 2 _GENERATED_85 _GENERATED_84 39 43 sram_filler $T=2014 -1150 0 0 $X=2018 $Y=-1150
XXB19A871F973 5 6 _GENERATED_87 _GENERATED_86 39 45 sram_filler $T=2466 -1024 0 180 $X=2018 $Y=-1613
XXB19A871F974 5 6 _GENERATED_89 _GENERATED_88 39 45 sram_filler $T=2802 -1024 0 180 $X=2354 $Y=-1613
XXB19A871F975 5 2 _GENERATED_91 _GENERATED_90 39 43 sram_filler $T=2350 -1150 0 0 $X=2354 $Y=-1150
XXB19A871F976 10 4 _GENERATED_93 _GENERATED_92 40 44 sram_filler $T=1794 824 0 180 $X=1346 $Y=234
XXB19A871F977 10 4 _GENERATED_95 _GENERATED_94 40 44 sram_filler $T=1458 824 0 180 $X=1010 $Y=234
XXB19A871F978 10 4 _GENERATED_97 _GENERATED_96 40 44 sram_filler $T=1122 824 0 180 $X=674 $Y=234
XXB19A871F979 10 4 _GENERATED_99 _GENERATED_98 40 44 sram_filler $T=786 824 0 180 $X=338 $Y=234
XXB19A871F980 10 4 _GENERATED_101 _GENERATED_100 40 44 sram_filler $T=450 824 0 180 $X=2 $Y=234
XXB19A871F981 10 7 7 _GENERATED_102 40 46 sram_filler $T=1342 698 0 0 $X=1346 $Y=698
XXB19A871F982 10 7 _GENERATED_103 10 40 46 sram_filler $T=1174 698 0 0 $X=1178 $Y=698
XXB19A871F983 10 7 _GENERATED_105 _GENERATED_104 40 46 sram_filler $T=838 698 0 0 $X=842 $Y=698
XXB19A871F984 10 7 7 _GENERATED_106 40 46 sram_filler $T=502 698 0 0 $X=506 $Y=698
XXB19A871F985 10 7 _GENERATED_107 10 40 46 sram_filler $T=334 698 0 0 $X=338 $Y=698
XXB19A871F986 10 7 _GENERATED_109 _GENERATED_108 40 46 sram_filler $T=-2 698 0 0 $X=2 $Y=698
XXB19A871F987 3 2 _GENERATED_110 3 41 43 sram_filler $T=2802 -100 0 180 $X=2354 $Y=-690
XXB19A871F988 3 2 2 _GENERATED_111 41 43 sram_filler $T=2634 -100 0 180 $X=2186 $Y=-690
XXB19A871F989 3 4 _GENERATED_112 3 41 44 sram_filler $T=2182 -226 0 0 $X=2186 $Y=-226
XXB19A871F990 3 4 4 _GENERATED_113 41 44 sram_filler $T=2350 -226 0 0 $X=2354 $Y=-226
XXB19A871F991 10 4 _GENERATED_114 10 40 44 sram_filler $T=2802 824 0 180 $X=2354 $Y=234
XXB19A871F992 10 4 4 _GENERATED_115 40 44 sram_filler $T=2634 824 0 180 $X=2186 $Y=234
XXB19A871F993 8 7 _GENERATED_116 8 42 46 sram_filler $T=2802 1748 0 180 $X=2354 $Y=1158
XXB19A871F994 8 7 7 _GENERATED_117 42 46 sram_filler $T=2634 1748 0 180 $X=2186 $Y=1158
XXB19A871F995 8 9 9 _GENERATED_118 42 47 sram_filler $T=2350 1622 0 0 $X=2354 $Y=1622
XXB19A871F996 8 9 _GENERATED_119 8 42 47 sram_filler $T=2182 1622 0 0 $X=2186 $Y=1622
XXB19A871F997 10 7 _GENERATED_120 10 40 46 sram_filler $T=1678 698 0 0 $X=1682 $Y=698
XXB19A871F998 10 4 4 _GENERATED_121 40 44 sram_filler $T=2130 824 0 180 $X=1682 $Y=234
.ends agen_unit
.subckt Write_Driver 2 3 4 6 7 8 9 10 11 12 13
+	14 15 16 17 18 19 20 21 22 23 24
+	25
MM1 3 25 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2386 $Y=852  $PIN_XY=2416,936,2386,852,2356,936 $DEVICE_ID=1001
MM2 10 25 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2218 $Y=852  $PIN_XY=2248,936,2218,852,2188,936 $DEVICE_ID=1001
MM3 3 8 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1546 $Y=1293  $PIN_XY=1576,1230,1546,1293,1516,1230 $DEVICE_ID=1001
MM4 3 7 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1546 $Y=873  $PIN_XY=1576,936,1546,873,1516,936 $DEVICE_ID=1001
MM5 9 8 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1378 $Y=1293  $PIN_XY=1408,1230,1378,1293,1348,1230 $DEVICE_ID=1001
MM6 25 7 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1378 $Y=852  $PIN_XY=1408,936,1378,852,1348,936 $DEVICE_ID=1001
MM7 8 12 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=874 $Y=1293  $PIN_XY=904,1230,874,1293,844,1230 $DEVICE_ID=1001
MM8 7 11 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=874 $Y=852  $PIN_XY=904,936,874,852,844,936 $DEVICE_ID=1001
MM9 12 6 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=370 $Y=1293  $PIN_XY=400,1230,370,1293,340,1230 $DEVICE_ID=1001
MM10 11 6 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=370 $Y=852  $PIN_XY=400,936,370,852,340,936 $DEVICE_ID=1001
XXB19A871F1031 2 3 10 25 7 21 22 23 buffer_highdrive $T=1154 1144 1 0 $X=1156 $Y=556
XXB19A871F1032 3 2 11 7 6 22 23 buffer $T=68 1148 1 0 $X=148 $Y=556
XXB19A871F1033 3 4 12 8 6 22 24 buffer $T=68 1018 0 0 $X=148 $Y=1020
XXB19A871F1034 3 2 17 18 22 23 sram_filler $T=3284 1146 0 180 $X=2836 $Y=556
XXB19A871F1035 3 4 19 20 22 24 sram_filler $T=3284 1020 1 180 $X=2836 $Y=1020
XXB19A871F1036 3 4 _GENERATED_26 5 22 24 sram_filler $T=2948 1020 1 180 $X=2500 $Y=1020
XXB19A871F1037 3 4 _GENERATED_27 5 22 24 sram_filler $T=2328 1020 0 0 $X=2332 $Y=1020
XXB19A871F1038 3 4 _GENERATED_29 _GENERATED_28 22 24 sram_filler $T=1992 1020 0 0 $X=1996 $Y=1020
XXB19A871F1039 3 4 9 8 22 24 invx4 $T=1132 1020 0 0 $X=1156 $Y=1020
.ends Write_Driver

* Hierarchy Level 0

* Top of hierarchy  cell=memory_array_static_column_decoder_test
.subckt memory_array_static_column_decoder_test GND! VDD! Q<1> Q<0> Q<2> Q<3> 8 9 10 11 12
+	13 14 15 16 17 18 19 20 21 22 23
+	24 25 26 27 28 29 30 31 32 33 34
+	35 36 37 38 39 73 74 75 76 77 78
+	79 80 81 82 83 84 85 86 87 88 89
+	90 91 92 93 94 95 96 97 98 WENB 100
+	101 102 103 104 WS0BAR 106 107 108 109 110 111
+	112 113 114 115 116 117 A<3> 119 120 121 122
+	123 124 CLK D<0> D<1> D<2> D<3> A<4> A<1> A<0> A<2>
MM1 GND! 460 273 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=14616  $PIN_XY=18174,14700,18144,14616,18114,14700 $DEVICE_ID=1001
MM2 38 124 460 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=14067  $PIN_XY=18174,14070,18144,14067,18114,14070 $DEVICE_ID=1001
MM3 GND! 458 268 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=13692  $PIN_XY=18174,13776,18144,13692,18114,13776 $DEVICE_ID=1001
MM4 38 123 458 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=13143  $PIN_XY=18174,13146,18144,13143,18114,13146 $DEVICE_ID=1001
MM5 GND! 453 262 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=12768  $PIN_XY=18174,12852,18144,12768,18114,12852 $DEVICE_ID=1001
MM6 38 122 453 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=12219  $PIN_XY=18174,12222,18144,12219,18114,12222 $DEVICE_ID=1001
MM7 GND! 411 259 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=11844  $PIN_XY=18174,11928,18144,11844,18114,11928 $DEVICE_ID=1001
MM8 273 124 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=14703  $PIN_XY=18006,14700,17976,14703,17946,14700 $DEVICE_ID=1001
MM9 460 273 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=14154  $PIN_XY=18006,14070,17976,14154,17946,14070 $DEVICE_ID=1001
MM10 268 123 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=13779  $PIN_XY=18006,13776,17976,13779,17946,13776 $DEVICE_ID=1001
MM11 458 268 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=13230  $PIN_XY=18006,13146,17976,13230,17946,13146 $DEVICE_ID=1001
MM12 262 122 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=12855  $PIN_XY=18006,12852,17976,12855,17946,12852 $DEVICE_ID=1001
MM13 453 262 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=12306  $PIN_XY=18006,12222,17976,12306,17946,12222 $DEVICE_ID=1001
MM14 259 121 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=11931  $PIN_XY=18006,11928,17976,11931,17946,11928 $DEVICE_ID=1001
MM15 GND! 461 272 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=14616  $PIN_XY=17502,14700,17472,14616,17442,14700 $DEVICE_ID=1001
MM16 36 124 461 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=14067  $PIN_XY=17502,14070,17472,14067,17442,14070 $DEVICE_ID=1001
MM17 GND! 457 267 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=13692  $PIN_XY=17502,13776,17472,13692,17442,13776 $DEVICE_ID=1001
MM18 36 123 457 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=13143  $PIN_XY=17502,13146,17472,13143,17442,13146 $DEVICE_ID=1001
MM19 GND! 452 263 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=12768  $PIN_XY=17502,12852,17472,12768,17442,12852 $DEVICE_ID=1001
MM20 36 122 452 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=12219  $PIN_XY=17502,12222,17472,12219,17442,12222 $DEVICE_ID=1001
MM21 GND! 412 260 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=11844  $PIN_XY=17502,11928,17472,11844,17442,11928 $DEVICE_ID=1001
MM22 272 124 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=14703  $PIN_XY=17334,14700,17304,14703,17274,14700 $DEVICE_ID=1001
MM23 461 272 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=14154  $PIN_XY=17334,14070,17304,14154,17274,14070 $DEVICE_ID=1001
MM24 267 123 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=13779  $PIN_XY=17334,13776,17304,13779,17274,13776 $DEVICE_ID=1001
MM25 457 267 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=13230  $PIN_XY=17334,13146,17304,13230,17274,13146 $DEVICE_ID=1001
MM26 263 122 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=12855  $PIN_XY=17334,12852,17304,12855,17274,12852 $DEVICE_ID=1001
MM27 452 263 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=12306  $PIN_XY=17334,12222,17304,12306,17274,12222 $DEVICE_ID=1001
MM28 260 121 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=11931  $PIN_XY=17334,11928,17304,11931,17274,11928 $DEVICE_ID=1001
MM29 GND! 462 271 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=14616  $PIN_XY=16830,14700,16800,14616,16770,14700 $DEVICE_ID=1001
MM30 34 124 462 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=14067  $PIN_XY=16830,14070,16800,14067,16770,14070 $DEVICE_ID=1001
MM31 GND! 456 266 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=13692  $PIN_XY=16830,13776,16800,13692,16770,13776 $DEVICE_ID=1001
MM32 34 123 456 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=13143  $PIN_XY=16830,13146,16800,13143,16770,13146 $DEVICE_ID=1001
MM33 GND! 451 264 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=12768  $PIN_XY=16830,12852,16800,12768,16770,12852 $DEVICE_ID=1001
MM34 34 122 451 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=12219  $PIN_XY=16830,12222,16800,12219,16770,12222 $DEVICE_ID=1001
MM35 GND! 413 261 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=11844  $PIN_XY=16830,11928,16800,11844,16770,11928 $DEVICE_ID=1001
MM36 271 124 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=14703  $PIN_XY=16662,14700,16632,14703,16602,14700 $DEVICE_ID=1001
MM37 462 271 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=14154  $PIN_XY=16662,14070,16632,14154,16602,14070 $DEVICE_ID=1001
MM38 266 123 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=13779  $PIN_XY=16662,13776,16632,13779,16602,13776 $DEVICE_ID=1001
MM39 456 266 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=13230  $PIN_XY=16662,13146,16632,13230,16602,13146 $DEVICE_ID=1001
MM40 264 122 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=12855  $PIN_XY=16662,12852,16632,12855,16602,12852 $DEVICE_ID=1001
MM41 451 264 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=12306  $PIN_XY=16662,12222,16632,12306,16602,12222 $DEVICE_ID=1001
MM42 261 121 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=11931  $PIN_XY=16662,11928,16632,11931,16602,11928 $DEVICE_ID=1001
MM43 38 121 411 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=11295  $PIN_XY=18174,11298,18144,11295,18114,11298 $DEVICE_ID=1001
MM44 GND! 408 257 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=10920  $PIN_XY=18174,11004,18144,10920,18114,11004 $DEVICE_ID=1001
MM45 38 120 408 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=10371  $PIN_XY=18174,10374,18144,10371,18114,10374 $DEVICE_ID=1001
MM46 GND! 406 187 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=9996  $PIN_XY=18174,10080,18144,9996,18114,10080 $DEVICE_ID=1001
MM47 38 119 406 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=9447  $PIN_XY=18174,9450,18144,9447,18114,9450 $DEVICE_ID=1001
MM48 GND! 363 186 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=9072  $PIN_XY=18174,9156,18144,9072,18114,9156 $DEVICE_ID=1001
MM49 38 116 363 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=8523  $PIN_XY=18174,8526,18144,8523,18114,8526 $DEVICE_ID=1001
MM50 411 259 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=11382  $PIN_XY=18006,11298,17976,11382,17946,11298 $DEVICE_ID=1001
MM51 257 120 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=11007  $PIN_XY=18006,11004,17976,11007,17946,11004 $DEVICE_ID=1001
MM52 408 257 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=10458  $PIN_XY=18006,10374,17976,10458,17946,10374 $DEVICE_ID=1001
MM53 187 119 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=10083  $PIN_XY=18006,10080,17976,10083,17946,10080 $DEVICE_ID=1001
MM54 406 187 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=9534  $PIN_XY=18006,9450,17976,9534,17946,9450 $DEVICE_ID=1001
MM55 186 116 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=9159  $PIN_XY=18006,9156,17976,9159,17946,9156 $DEVICE_ID=1001
MM56 363 186 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=8610  $PIN_XY=18006,8526,17976,8610,17946,8526 $DEVICE_ID=1001
MM57 36 121 412 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=11295  $PIN_XY=17502,11298,17472,11295,17442,11298 $DEVICE_ID=1001
MM58 GND! 409 256 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=10920  $PIN_XY=17502,11004,17472,10920,17442,11004 $DEVICE_ID=1001
MM59 36 120 409 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=10371  $PIN_XY=17502,10374,17472,10371,17442,10374 $DEVICE_ID=1001
MM60 GND! 405 189 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=9996  $PIN_XY=17502,10080,17472,9996,17442,10080 $DEVICE_ID=1001
MM61 36 119 405 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=9447  $PIN_XY=17502,9450,17472,9447,17442,9450 $DEVICE_ID=1001
MM62 GND! 364 188 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=9072  $PIN_XY=17502,9156,17472,9072,17442,9156 $DEVICE_ID=1001
MM63 36 116 364 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=8523  $PIN_XY=17502,8526,17472,8523,17442,8526 $DEVICE_ID=1001
MM64 412 260 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=11382  $PIN_XY=17334,11298,17304,11382,17274,11298 $DEVICE_ID=1001
MM65 256 120 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=11007  $PIN_XY=17334,11004,17304,11007,17274,11004 $DEVICE_ID=1001
MM66 409 256 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=10458  $PIN_XY=17334,10374,17304,10458,17274,10374 $DEVICE_ID=1001
MM67 189 119 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=10083  $PIN_XY=17334,10080,17304,10083,17274,10080 $DEVICE_ID=1001
MM68 405 189 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=9534  $PIN_XY=17334,9450,17304,9534,17274,9450 $DEVICE_ID=1001
MM69 188 116 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=9159  $PIN_XY=17334,9156,17304,9159,17274,9156 $DEVICE_ID=1001
MM70 364 188 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=8610  $PIN_XY=17334,8526,17304,8610,17274,8526 $DEVICE_ID=1001
MM71 34 121 413 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=11295  $PIN_XY=16830,11298,16800,11295,16770,11298 $DEVICE_ID=1001
MM72 GND! 410 255 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=10920  $PIN_XY=16830,11004,16800,10920,16770,11004 $DEVICE_ID=1001
MM73 34 120 410 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=10371  $PIN_XY=16830,10374,16800,10371,16770,10374 $DEVICE_ID=1001
MM74 GND! 404 191 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=9996  $PIN_XY=16830,10080,16800,9996,16770,10080 $DEVICE_ID=1001
MM75 34 119 404 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=9447  $PIN_XY=16830,9450,16800,9447,16770,9450 $DEVICE_ID=1001
MM76 GND! 365 190 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=9072  $PIN_XY=16830,9156,16800,9072,16770,9156 $DEVICE_ID=1001
MM77 34 116 365 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=8523  $PIN_XY=16830,8526,16800,8523,16770,8526 $DEVICE_ID=1001
MM78 413 261 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=11382  $PIN_XY=16662,11298,16632,11382,16602,11298 $DEVICE_ID=1001
MM79 255 120 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=11007  $PIN_XY=16662,11004,16632,11007,16602,11004 $DEVICE_ID=1001
MM80 410 255 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=10458  $PIN_XY=16662,10374,16632,10458,16602,10374 $DEVICE_ID=1001
MM81 191 119 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=10083  $PIN_XY=16662,10080,16632,10083,16602,10080 $DEVICE_ID=1001
MM82 404 191 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=9534  $PIN_XY=16662,9450,16632,9534,16602,9450 $DEVICE_ID=1001
MM83 190 116 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=9159  $PIN_XY=16662,9156,16632,9159,16602,9156 $DEVICE_ID=1001
MM84 365 190 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=8610  $PIN_XY=16662,8526,16632,8610,16602,8526 $DEVICE_ID=1001
MM85 GND! 459 270 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=14616  $PIN_XY=16158,14700,16128,14616,16098,14700 $DEVICE_ID=1001
MM86 32 124 459 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=14067  $PIN_XY=16158,14070,16128,14067,16098,14070 $DEVICE_ID=1001
MM87 GND! 455 269 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=13692  $PIN_XY=16158,13776,16128,13692,16098,13776 $DEVICE_ID=1001
MM88 32 123 455 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=13143  $PIN_XY=16158,13146,16128,13143,16098,13146 $DEVICE_ID=1001
MM89 GND! 454 265 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=12768  $PIN_XY=16158,12852,16128,12768,16098,12852 $DEVICE_ID=1001
MM90 32 122 454 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=12219  $PIN_XY=16158,12222,16128,12219,16098,12222 $DEVICE_ID=1001
MM91 GND! 414 258 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=11844  $PIN_XY=16158,11928,16128,11844,16098,11928 $DEVICE_ID=1001
MM92 270 124 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=14703  $PIN_XY=15990,14700,15960,14703,15930,14700 $DEVICE_ID=1001
MM93 459 270 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=14154  $PIN_XY=15990,14070,15960,14154,15930,14070 $DEVICE_ID=1001
MM94 269 123 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=13779  $PIN_XY=15990,13776,15960,13779,15930,13776 $DEVICE_ID=1001
MM95 455 269 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=13230  $PIN_XY=15990,13146,15960,13230,15930,13146 $DEVICE_ID=1001
MM96 265 122 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=12855  $PIN_XY=15990,12852,15960,12855,15930,12852 $DEVICE_ID=1001
MM97 454 265 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=12306  $PIN_XY=15990,12222,15960,12306,15930,12222 $DEVICE_ID=1001
MM98 258 121 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=11931  $PIN_XY=15990,11928,15960,11931,15930,11928 $DEVICE_ID=1001
MM99 GND! 463 234 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=14616  $PIN_XY=15150,14700,15120,14616,15090,14700 $DEVICE_ID=1001
MM100 31 124 463 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=14067  $PIN_XY=15150,14070,15120,14067,15090,14070 $DEVICE_ID=1001
MM101 GND! 464 235 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=13692  $PIN_XY=15150,13776,15120,13692,15090,13776 $DEVICE_ID=1001
MM102 31 123 464 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=13143  $PIN_XY=15150,13146,15120,13143,15090,13146 $DEVICE_ID=1001
MM103 GND! 465 236 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=12768  $PIN_XY=15150,12852,15120,12768,15090,12852 $DEVICE_ID=1001
MM104 31 122 465 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=12219  $PIN_XY=15150,12222,15120,12219,15090,12222 $DEVICE_ID=1001
MM105 GND! 415 237 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=11844  $PIN_XY=15150,11928,15120,11844,15090,11928 $DEVICE_ID=1001
MM106 234 124 30 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=14703  $PIN_XY=14982,14700,14952,14703,14922,14700 $DEVICE_ID=1001
MM107 463 234 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=14154  $PIN_XY=14982,14070,14952,14154,14922,14070 $DEVICE_ID=1001
MM108 235 123 30 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=13779  $PIN_XY=14982,13776,14952,13779,14922,13776 $DEVICE_ID=1001
MM109 464 235 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=13230  $PIN_XY=14982,13146,14952,13230,14922,13146 $DEVICE_ID=1001
MM110 236 122 30 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=12855  $PIN_XY=14982,12852,14952,12855,14922,12852 $DEVICE_ID=1001
MM111 465 236 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=12306  $PIN_XY=14982,12222,14952,12306,14922,12222 $DEVICE_ID=1001
MM112 237 121 30 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=11931  $PIN_XY=14982,11928,14952,11931,14922,11928 $DEVICE_ID=1001
MM113 GND! 467 240 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=14616  $PIN_XY=14478,14700,14448,14616,14418,14700 $DEVICE_ID=1001
MM114 24 124 467 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=14067  $PIN_XY=14478,14070,14448,14067,14418,14070 $DEVICE_ID=1001
MM115 GND! 469 242 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=13692  $PIN_XY=14478,13776,14448,13692,14418,13776 $DEVICE_ID=1001
MM116 24 123 469 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=13143  $PIN_XY=14478,13146,14448,13143,14418,13146 $DEVICE_ID=1001
MM117 GND! 473 246 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=12768  $PIN_XY=14478,12852,14448,12768,14418,12852 $DEVICE_ID=1001
MM118 24 122 473 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=12219  $PIN_XY=14478,12222,14448,12219,14418,12222 $DEVICE_ID=1001
MM119 GND! 420 250 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=11844  $PIN_XY=14478,11928,14448,11844,14418,11928 $DEVICE_ID=1001
MM120 240 124 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=14703  $PIN_XY=14310,14700,14280,14703,14250,14700 $DEVICE_ID=1001
MM121 467 240 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=14154  $PIN_XY=14310,14070,14280,14154,14250,14070 $DEVICE_ID=1001
MM122 242 123 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=13779  $PIN_XY=14310,13776,14280,13779,14250,13776 $DEVICE_ID=1001
MM123 469 242 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=13230  $PIN_XY=14310,13146,14280,13230,14250,13146 $DEVICE_ID=1001
MM124 246 122 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=12855  $PIN_XY=14310,12852,14280,12855,14250,12852 $DEVICE_ID=1001
MM125 473 246 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=12306  $PIN_XY=14310,12222,14280,12306,14250,12222 $DEVICE_ID=1001
MM126 250 121 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=11931  $PIN_XY=14310,11928,14280,11931,14250,11928 $DEVICE_ID=1001
MM127 32 121 414 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=11295  $PIN_XY=16158,11298,16128,11295,16098,11298 $DEVICE_ID=1001
MM128 GND! 407 254 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=10920  $PIN_XY=16158,11004,16128,10920,16098,11004 $DEVICE_ID=1001
MM129 32 120 407 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=10371  $PIN_XY=16158,10374,16128,10371,16098,10374 $DEVICE_ID=1001
MM130 GND! 403 193 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=9996  $PIN_XY=16158,10080,16128,9996,16098,10080 $DEVICE_ID=1001
MM131 32 119 403 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=9447  $PIN_XY=16158,9450,16128,9447,16098,9450 $DEVICE_ID=1001
MM132 GND! 366 192 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=9072  $PIN_XY=16158,9156,16128,9072,16098,9156 $DEVICE_ID=1001
MM133 32 116 366 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=8523  $PIN_XY=16158,8526,16128,8523,16098,8526 $DEVICE_ID=1001
MM134 414 258 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=11382  $PIN_XY=15990,11298,15960,11382,15930,11298 $DEVICE_ID=1001
MM135 254 120 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=11007  $PIN_XY=15990,11004,15960,11007,15930,11004 $DEVICE_ID=1001
MM136 407 254 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=10458  $PIN_XY=15990,10374,15960,10458,15930,10374 $DEVICE_ID=1001
MM137 193 119 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=10083  $PIN_XY=15990,10080,15960,10083,15930,10080 $DEVICE_ID=1001
MM138 403 193 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=9534  $PIN_XY=15990,9450,15960,9534,15930,9450 $DEVICE_ID=1001
MM139 192 116 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=9159  $PIN_XY=15990,9156,15960,9159,15930,9156 $DEVICE_ID=1001
MM140 366 192 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=8610  $PIN_XY=15990,8526,15960,8610,15930,8526 $DEVICE_ID=1001
MM141 31 121 415 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=11295  $PIN_XY=15150,11298,15120,11295,15090,11298 $DEVICE_ID=1001
MM142 GND! 416 238 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=10920  $PIN_XY=15150,11004,15120,10920,15090,11004 $DEVICE_ID=1001
MM143 31 120 416 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=10371  $PIN_XY=15150,10374,15120,10371,15090,10374 $DEVICE_ID=1001
MM144 GND! 417 175 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=9996  $PIN_XY=15150,10080,15120,9996,15090,10080 $DEVICE_ID=1001
MM145 31 119 417 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=9447  $PIN_XY=15150,9450,15120,9447,15090,9450 $DEVICE_ID=1001
MM146 GND! 367 174 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=9072  $PIN_XY=15150,9156,15120,9072,15090,9156 $DEVICE_ID=1001
MM147 31 116 367 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=8523  $PIN_XY=15150,8526,15120,8523,15090,8526 $DEVICE_ID=1001
MM148 415 237 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=11382  $PIN_XY=14982,11298,14952,11382,14922,11298 $DEVICE_ID=1001
MM149 238 120 30 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=11007  $PIN_XY=14982,11004,14952,11007,14922,11004 $DEVICE_ID=1001
MM150 416 238 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=10458  $PIN_XY=14982,10374,14952,10458,14922,10374 $DEVICE_ID=1001
MM151 175 119 30 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=10083  $PIN_XY=14982,10080,14952,10083,14922,10080 $DEVICE_ID=1001
MM152 417 175 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=9534  $PIN_XY=14982,9450,14952,9534,14922,9450 $DEVICE_ID=1001
MM153 174 116 30 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=9159  $PIN_XY=14982,9156,14952,9159,14922,9156 $DEVICE_ID=1001
MM154 367 174 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=8610  $PIN_XY=14982,8526,14952,8610,14922,8526 $DEVICE_ID=1001
MM155 24 121 420 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=11295  $PIN_XY=14478,11298,14448,11295,14418,11298 $DEVICE_ID=1001
MM156 GND! 422 252 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=10920  $PIN_XY=14478,11004,14448,10920,14418,11004 $DEVICE_ID=1001
MM157 24 120 422 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=10371  $PIN_XY=14478,10374,14448,10371,14418,10374 $DEVICE_ID=1001
MM158 GND! 424 181 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=9996  $PIN_XY=14478,10080,14448,9996,14418,10080 $DEVICE_ID=1001
MM159 24 119 424 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=9447  $PIN_XY=14478,9450,14448,9447,14418,9450 $DEVICE_ID=1001
MM160 GND! 374 180 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=9072  $PIN_XY=14478,9156,14448,9072,14418,9156 $DEVICE_ID=1001
MM161 24 116 374 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=8523  $PIN_XY=14478,8526,14448,8523,14418,8526 $DEVICE_ID=1001
MM162 420 250 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=11382  $PIN_XY=14310,11298,14280,11382,14250,11298 $DEVICE_ID=1001
MM163 252 120 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=11007  $PIN_XY=14310,11004,14280,11007,14250,11004 $DEVICE_ID=1001
MM164 422 252 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=10458  $PIN_XY=14310,10374,14280,10458,14250,10374 $DEVICE_ID=1001
MM165 181 119 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=10083  $PIN_XY=14310,10080,14280,10083,14250,10080 $DEVICE_ID=1001
MM166 424 181 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=9534  $PIN_XY=14310,9450,14280,9534,14250,9450 $DEVICE_ID=1001
MM167 180 116 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=9159  $PIN_XY=14310,9156,14280,9159,14250,9156 $DEVICE_ID=1001
MM168 374 180 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=8610  $PIN_XY=14310,8526,14280,8610,14250,8526 $DEVICE_ID=1001
MM169 GND! 466 239 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=14616  $PIN_XY=13806,14700,13776,14616,13746,14700 $DEVICE_ID=1001
MM170 26 124 466 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=14067  $PIN_XY=13806,14070,13776,14067,13746,14070 $DEVICE_ID=1001
MM171 GND! 470 243 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=13692  $PIN_XY=13806,13776,13776,13692,13746,13776 $DEVICE_ID=1001
MM172 26 123 470 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=13143  $PIN_XY=13806,13146,13776,13143,13746,13146 $DEVICE_ID=1001
MM173 GND! 474 247 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=12768  $PIN_XY=13806,12852,13776,12768,13746,12852 $DEVICE_ID=1001
MM174 26 122 474 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=12219  $PIN_XY=13806,12222,13776,12219,13746,12222 $DEVICE_ID=1001
MM175 GND! 419 249 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=11844  $PIN_XY=13806,11928,13776,11844,13746,11928 $DEVICE_ID=1001
MM176 26 121 419 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=11295  $PIN_XY=13806,11298,13776,11295,13746,11298 $DEVICE_ID=1001
MM177 GND! 421 251 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=10920  $PIN_XY=13806,11004,13776,10920,13746,11004 $DEVICE_ID=1001
MM178 26 120 421 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=10371  $PIN_XY=13806,10374,13776,10371,13746,10374 $DEVICE_ID=1001
MM179 GND! 425 179 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=9996  $PIN_XY=13806,10080,13776,9996,13746,10080 $DEVICE_ID=1001
MM180 26 119 425 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=9447  $PIN_XY=13806,9450,13776,9447,13746,9450 $DEVICE_ID=1001
MM181 GND! 373 178 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=9072  $PIN_XY=13806,9156,13776,9072,13746,9156 $DEVICE_ID=1001
MM182 26 116 373 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=8523  $PIN_XY=13806,8526,13776,8523,13746,8526 $DEVICE_ID=1001
MM183 239 124 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=14703  $PIN_XY=13638,14700,13608,14703,13578,14700 $DEVICE_ID=1001
MM184 466 239 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=14154  $PIN_XY=13638,14070,13608,14154,13578,14070 $DEVICE_ID=1001
MM185 243 123 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=13779  $PIN_XY=13638,13776,13608,13779,13578,13776 $DEVICE_ID=1001
MM186 470 243 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=13230  $PIN_XY=13638,13146,13608,13230,13578,13146 $DEVICE_ID=1001
MM187 247 122 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=12855  $PIN_XY=13638,12852,13608,12855,13578,12852 $DEVICE_ID=1001
MM188 474 247 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=12306  $PIN_XY=13638,12222,13608,12306,13578,12222 $DEVICE_ID=1001
MM189 249 121 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=11931  $PIN_XY=13638,11928,13608,11931,13578,11928 $DEVICE_ID=1001
MM190 419 249 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=11382  $PIN_XY=13638,11298,13608,11382,13578,11298 $DEVICE_ID=1001
MM191 251 120 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=11007  $PIN_XY=13638,11004,13608,11007,13578,11004 $DEVICE_ID=1001
MM192 421 251 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=10458  $PIN_XY=13638,10374,13608,10458,13578,10374 $DEVICE_ID=1001
MM193 179 119 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=10083  $PIN_XY=13638,10080,13608,10083,13578,10080 $DEVICE_ID=1001
MM194 425 179 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=9534  $PIN_XY=13638,9450,13608,9534,13578,9450 $DEVICE_ID=1001
MM195 178 116 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=9159  $PIN_XY=13638,9156,13608,9159,13578,9156 $DEVICE_ID=1001
MM196 373 178 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=8610  $PIN_XY=13638,8526,13608,8610,13578,8526 $DEVICE_ID=1001
MM197 GND! 468 241 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=14616  $PIN_XY=13134,14700,13104,14616,13074,14700 $DEVICE_ID=1001
MM198 28 124 468 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=14067  $PIN_XY=13134,14070,13104,14067,13074,14070 $DEVICE_ID=1001
MM199 GND! 471 244 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=13692  $PIN_XY=13134,13776,13104,13692,13074,13776 $DEVICE_ID=1001
MM200 28 123 471 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=13143  $PIN_XY=13134,13146,13104,13143,13074,13146 $DEVICE_ID=1001
MM201 GND! 472 245 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=12768  $PIN_XY=13134,12852,13104,12768,13074,12852 $DEVICE_ID=1001
MM202 28 122 472 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=12219  $PIN_XY=13134,12222,13104,12219,13074,12222 $DEVICE_ID=1001
MM203 GND! 418 248 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=11844  $PIN_XY=13134,11928,13104,11844,13074,11928 $DEVICE_ID=1001
MM204 28 121 418 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=11295  $PIN_XY=13134,11298,13104,11295,13074,11298 $DEVICE_ID=1001
MM205 GND! 423 253 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=10920  $PIN_XY=13134,11004,13104,10920,13074,11004 $DEVICE_ID=1001
MM206 28 120 423 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=10371  $PIN_XY=13134,10374,13104,10371,13074,10374 $DEVICE_ID=1001
MM207 GND! 426 177 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=9996  $PIN_XY=13134,10080,13104,9996,13074,10080 $DEVICE_ID=1001
MM208 28 119 426 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=9447  $PIN_XY=13134,9450,13104,9447,13074,9450 $DEVICE_ID=1001
MM209 GND! 372 176 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=9072  $PIN_XY=13134,9156,13104,9072,13074,9156 $DEVICE_ID=1001
MM210 28 116 372 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=8523  $PIN_XY=13134,8526,13104,8523,13074,8526 $DEVICE_ID=1001
MM211 241 124 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=14703  $PIN_XY=12966,14700,12936,14703,12906,14700 $DEVICE_ID=1001
MM212 468 241 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=14154  $PIN_XY=12966,14070,12936,14154,12906,14070 $DEVICE_ID=1001
MM213 244 123 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=13779  $PIN_XY=12966,13776,12936,13779,12906,13776 $DEVICE_ID=1001
MM214 471 244 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=13230  $PIN_XY=12966,13146,12936,13230,12906,13146 $DEVICE_ID=1001
MM215 245 122 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=12855  $PIN_XY=12966,12852,12936,12855,12906,12852 $DEVICE_ID=1001
MM216 472 245 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=12306  $PIN_XY=12966,12222,12936,12306,12906,12222 $DEVICE_ID=1001
MM217 248 121 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=11931  $PIN_XY=12966,11928,12936,11931,12906,11928 $DEVICE_ID=1001
MM218 418 248 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=11382  $PIN_XY=12966,11298,12936,11382,12906,11298 $DEVICE_ID=1001
MM219 253 120 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=11007  $PIN_XY=12966,11004,12936,11007,12906,11004 $DEVICE_ID=1001
MM220 423 253 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=10458  $PIN_XY=12966,10374,12936,10458,12906,10374 $DEVICE_ID=1001
MM221 177 119 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=10083  $PIN_XY=12966,10080,12936,10083,12906,10080 $DEVICE_ID=1001
MM222 426 177 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=9534  $PIN_XY=12966,9450,12936,9534,12906,9450 $DEVICE_ID=1001
MM223 176 116 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=9159  $PIN_XY=12966,9156,12936,9159,12906,9156 $DEVICE_ID=1001
MM224 372 176 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=8610  $PIN_XY=12966,8526,12936,8610,12906,8526 $DEVICE_ID=1001
MM225 GND! 441 216 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=14616  $PIN_XY=12126,14700,12096,14616,12066,14700 $DEVICE_ID=1001
MM226 23 124 441 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=14067  $PIN_XY=12126,14070,12096,14067,12066,14070 $DEVICE_ID=1001
MM227 GND! 443 218 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=13692  $PIN_XY=12126,13776,12096,13692,12066,13776 $DEVICE_ID=1001
MM228 23 123 443 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=13143  $PIN_XY=12126,13146,12096,13143,12066,13146 $DEVICE_ID=1001
MM229 GND! 448 223 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=12768  $PIN_XY=12126,12852,12096,12768,12066,12852 $DEVICE_ID=1001
MM230 23 122 448 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=12219  $PIN_XY=12126,12222,12096,12219,12066,12222 $DEVICE_ID=1001
MM231 GND! 394 229 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=11844  $PIN_XY=12126,11928,12096,11844,12066,11928 $DEVICE_ID=1001
MM232 216 124 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=14703  $PIN_XY=11958,14700,11928,14703,11898,14700 $DEVICE_ID=1001
MM233 441 216 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=14154  $PIN_XY=11958,14070,11928,14154,11898,14070 $DEVICE_ID=1001
MM234 218 123 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=13779  $PIN_XY=11958,13776,11928,13779,11898,13776 $DEVICE_ID=1001
MM235 443 218 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=13230  $PIN_XY=11958,13146,11928,13230,11898,13146 $DEVICE_ID=1001
MM236 223 122 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=12855  $PIN_XY=11958,12852,11928,12855,11898,12852 $DEVICE_ID=1001
MM237 448 223 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=12306  $PIN_XY=11958,12222,11928,12306,11898,12222 $DEVICE_ID=1001
MM238 229 121 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=11931  $PIN_XY=11958,11928,11928,11931,11898,11928 $DEVICE_ID=1001
MM239 GND! 440 215 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=14616  $PIN_XY=11454,14700,11424,14616,11394,14700 $DEVICE_ID=1001
MM240 21 124 440 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=14067  $PIN_XY=11454,14070,11424,14067,11394,14070 $DEVICE_ID=1001
MM241 GND! 444 219 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=13692  $PIN_XY=11454,13776,11424,13692,11394,13776 $DEVICE_ID=1001
MM242 21 123 444 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=13143  $PIN_XY=11454,13146,11424,13143,11394,13146 $DEVICE_ID=1001
MM243 GND! 449 224 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=12768  $PIN_XY=11454,12852,11424,12768,11394,12852 $DEVICE_ID=1001
MM244 21 122 449 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=12219  $PIN_XY=11454,12222,11424,12219,11394,12222 $DEVICE_ID=1001
MM245 GND! 393 228 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=11844  $PIN_XY=11454,11928,11424,11844,11394,11928 $DEVICE_ID=1001
MM246 215 124 20 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=14703  $PIN_XY=11286,14700,11256,14703,11226,14700 $DEVICE_ID=1001
MM247 440 215 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=14154  $PIN_XY=11286,14070,11256,14154,11226,14070 $DEVICE_ID=1001
MM248 219 123 20 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=13779  $PIN_XY=11286,13776,11256,13779,11226,13776 $DEVICE_ID=1001
MM249 444 219 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=13230  $PIN_XY=11286,13146,11256,13230,11226,13146 $DEVICE_ID=1001
MM250 224 122 20 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=12855  $PIN_XY=11286,12852,11256,12855,11226,12852 $DEVICE_ID=1001
MM251 449 224 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=12306  $PIN_XY=11286,12222,11256,12306,11226,12222 $DEVICE_ID=1001
MM252 228 121 20 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=11931  $PIN_XY=11286,11928,11256,11931,11226,11928 $DEVICE_ID=1001
MM253 GND! 439 214 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=14616  $PIN_XY=10782,14700,10752,14616,10722,14700 $DEVICE_ID=1001
MM254 19 124 439 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=14067  $PIN_XY=10782,14070,10752,14067,10722,14070 $DEVICE_ID=1001
MM255 GND! 445 220 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=13692  $PIN_XY=10782,13776,10752,13692,10722,13776 $DEVICE_ID=1001
MM256 19 123 445 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=13143  $PIN_XY=10782,13146,10752,13143,10722,13146 $DEVICE_ID=1001
MM257 GND! 450 225 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=12768  $PIN_XY=10782,12852,10752,12768,10722,12852 $DEVICE_ID=1001
MM258 19 122 450 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=12219  $PIN_XY=10782,12222,10752,12219,10722,12222 $DEVICE_ID=1001
MM259 GND! 392 227 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=11844  $PIN_XY=10782,11928,10752,11844,10722,11928 $DEVICE_ID=1001
MM260 214 124 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=14703  $PIN_XY=10614,14700,10584,14703,10554,14700 $DEVICE_ID=1001
MM261 439 214 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=14154  $PIN_XY=10614,14070,10584,14154,10554,14070 $DEVICE_ID=1001
MM262 220 123 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=13779  $PIN_XY=10614,13776,10584,13779,10554,13776 $DEVICE_ID=1001
MM263 445 220 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=13230  $PIN_XY=10614,13146,10584,13230,10554,13146 $DEVICE_ID=1001
MM264 225 122 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=12855  $PIN_XY=10614,12852,10584,12855,10554,12852 $DEVICE_ID=1001
MM265 450 225 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=12306  $PIN_XY=10614,12222,10584,12306,10554,12222 $DEVICE_ID=1001
MM266 227 121 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=11931  $PIN_XY=10614,11928,10584,11931,10554,11928 $DEVICE_ID=1001
MM267 23 121 394 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=11295  $PIN_XY=12126,11298,12096,11295,12066,11298 $DEVICE_ID=1001
MM268 GND! 397 232 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=10920  $PIN_XY=12126,11004,12096,10920,12066,11004 $DEVICE_ID=1001
MM269 23 120 397 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=10371  $PIN_XY=12126,10374,12096,10371,12066,10374 $DEVICE_ID=1001
MM270 GND! 399 169 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=9996  $PIN_XY=12126,10080,12096,9996,12066,10080 $DEVICE_ID=1001
MM271 23 119 399 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=9447  $PIN_XY=12126,9450,12096,9447,12066,9450 $DEVICE_ID=1001
MM272 GND! 358 168 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=9072  $PIN_XY=12126,9156,12096,9072,12066,9156 $DEVICE_ID=1001
MM273 23 116 358 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=8523  $PIN_XY=12126,8526,12096,8523,12066,8526 $DEVICE_ID=1001
MM274 394 229 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=11382  $PIN_XY=11958,11298,11928,11382,11898,11298 $DEVICE_ID=1001
MM275 232 120 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=11007  $PIN_XY=11958,11004,11928,11007,11898,11004 $DEVICE_ID=1001
MM276 397 232 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=10458  $PIN_XY=11958,10374,11928,10458,11898,10374 $DEVICE_ID=1001
MM277 169 119 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=10083  $PIN_XY=11958,10080,11928,10083,11898,10080 $DEVICE_ID=1001
MM278 399 169 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=9534  $PIN_XY=11958,9450,11928,9534,11898,9450 $DEVICE_ID=1001
MM279 168 116 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=9159  $PIN_XY=11958,9156,11928,9159,11898,9156 $DEVICE_ID=1001
MM280 358 168 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=8610  $PIN_XY=11958,8526,11928,8610,11898,8526 $DEVICE_ID=1001
MM281 21 121 393 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=11295  $PIN_XY=11454,11298,11424,11295,11394,11298 $DEVICE_ID=1001
MM282 GND! 396 231 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=10920  $PIN_XY=11454,11004,11424,10920,11394,11004 $DEVICE_ID=1001
MM283 21 120 396 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=10371  $PIN_XY=11454,10374,11424,10371,11394,10374 $DEVICE_ID=1001
MM284 GND! 400 167 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=9996  $PIN_XY=11454,10080,11424,9996,11394,10080 $DEVICE_ID=1001
MM285 21 119 400 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=9447  $PIN_XY=11454,9450,11424,9447,11394,9450 $DEVICE_ID=1001
MM286 GND! 357 166 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=9072  $PIN_XY=11454,9156,11424,9072,11394,9156 $DEVICE_ID=1001
MM287 21 116 357 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=8523  $PIN_XY=11454,8526,11424,8523,11394,8526 $DEVICE_ID=1001
MM288 393 228 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=11382  $PIN_XY=11286,11298,11256,11382,11226,11298 $DEVICE_ID=1001
MM289 231 120 20 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=11007  $PIN_XY=11286,11004,11256,11007,11226,11004 $DEVICE_ID=1001
MM290 396 231 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=10458  $PIN_XY=11286,10374,11256,10458,11226,10374 $DEVICE_ID=1001
MM291 167 119 20 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=10083  $PIN_XY=11286,10080,11256,10083,11226,10080 $DEVICE_ID=1001
MM292 400 167 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=9534  $PIN_XY=11286,9450,11256,9534,11226,9450 $DEVICE_ID=1001
MM293 166 116 20 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=9159  $PIN_XY=11286,9156,11256,9159,11226,9156 $DEVICE_ID=1001
MM294 357 166 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=8610  $PIN_XY=11286,8526,11256,8610,11226,8526 $DEVICE_ID=1001
MM295 19 121 392 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=11295  $PIN_XY=10782,11298,10752,11295,10722,11298 $DEVICE_ID=1001
MM296 GND! 395 230 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=10920  $PIN_XY=10782,11004,10752,10920,10722,11004 $DEVICE_ID=1001
MM297 19 120 395 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=10371  $PIN_XY=10782,10374,10752,10371,10722,10374 $DEVICE_ID=1001
MM298 GND! 401 165 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=9996  $PIN_XY=10782,10080,10752,9996,10722,10080 $DEVICE_ID=1001
MM299 19 119 401 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=9447  $PIN_XY=10782,9450,10752,9447,10722,9450 $DEVICE_ID=1001
MM300 GND! 356 164 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=9072  $PIN_XY=10782,9156,10752,9072,10722,9156 $DEVICE_ID=1001
MM301 19 116 356 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=8523  $PIN_XY=10782,8526,10752,8523,10722,8526 $DEVICE_ID=1001
MM302 392 227 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=11382  $PIN_XY=10614,11298,10584,11382,10554,11298 $DEVICE_ID=1001
MM303 230 120 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=11007  $PIN_XY=10614,11004,10584,11007,10554,11004 $DEVICE_ID=1001
MM304 395 230 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=10458  $PIN_XY=10614,10374,10584,10458,10554,10374 $DEVICE_ID=1001
MM305 165 119 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=10083  $PIN_XY=10614,10080,10584,10083,10554,10080 $DEVICE_ID=1001
MM306 401 165 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=9534  $PIN_XY=10614,9450,10584,9534,10554,9450 $DEVICE_ID=1001
MM307 164 116 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=9159  $PIN_XY=10614,9156,10584,9159,10554,9156 $DEVICE_ID=1001
MM308 356 164 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=8610  $PIN_XY=10614,8526,10584,8610,10554,8526 $DEVICE_ID=1001
MM309 GND! 442 217 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=14616  $PIN_XY=10110,14700,10080,14616,10050,14700 $DEVICE_ID=1001
MM310 16 124 442 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=14067  $PIN_XY=10110,14070,10080,14067,10050,14070 $DEVICE_ID=1001
MM311 GND! 446 221 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=13692  $PIN_XY=10110,13776,10080,13692,10050,13776 $DEVICE_ID=1001
MM312 16 123 446 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=13143  $PIN_XY=10110,13146,10080,13143,10050,13146 $DEVICE_ID=1001
MM313 GND! 447 222 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=12768  $PIN_XY=10110,12852,10080,12768,10050,12852 $DEVICE_ID=1001
MM314 16 122 447 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=12219  $PIN_XY=10110,12222,10080,12219,10050,12222 $DEVICE_ID=1001
MM315 GND! 391 226 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=11844  $PIN_XY=10110,11928,10080,11844,10050,11928 $DEVICE_ID=1001
MM316 217 124 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=14703  $PIN_XY=9942,14700,9912,14703,9882,14700 $DEVICE_ID=1001
MM317 442 217 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=14154  $PIN_XY=9942,14070,9912,14154,9882,14070 $DEVICE_ID=1001
MM318 221 123 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=13779  $PIN_XY=9942,13776,9912,13779,9882,13776 $DEVICE_ID=1001
MM319 446 221 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=13230  $PIN_XY=9942,13146,9912,13230,9882,13146 $DEVICE_ID=1001
MM320 222 122 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=12855  $PIN_XY=9942,12852,9912,12855,9882,12852 $DEVICE_ID=1001
MM321 447 222 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=12306  $PIN_XY=9942,12222,9912,12306,9882,12222 $DEVICE_ID=1001
MM322 226 121 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=11931  $PIN_XY=9942,11928,9912,11931,9882,11928 $DEVICE_ID=1001
MM323 GND! 436 213 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=14616  $PIN_XY=9102,14700,9072,14616,9042,14700 $DEVICE_ID=1001
MM324 8 124 436 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=14067  $PIN_XY=9102,14070,9072,14067,9042,14070 $DEVICE_ID=1001
MM325 GND! 434 208 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=13692  $PIN_XY=9102,13776,9072,13692,9042,13776 $DEVICE_ID=1001
MM326 8 123 434 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=13143  $PIN_XY=9102,13146,9072,13143,9042,13146 $DEVICE_ID=1001
MM327 GND! 429 202 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=12768  $PIN_XY=9102,12852,9072,12768,9042,12852 $DEVICE_ID=1001
MM328 8 122 429 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=12219  $PIN_XY=9102,12222,9072,12219,9042,12222 $DEVICE_ID=1001
MM329 GND! 387 199 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=11844  $PIN_XY=9102,11928,9072,11844,9042,11928 $DEVICE_ID=1001
MM330 213 124 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=14703  $PIN_XY=8934,14700,8904,14703,8874,14700 $DEVICE_ID=1001
MM331 436 213 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=14154  $PIN_XY=8934,14070,8904,14154,8874,14070 $DEVICE_ID=1001
MM332 208 123 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=13779  $PIN_XY=8934,13776,8904,13779,8874,13776 $DEVICE_ID=1001
MM333 434 208 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=13230  $PIN_XY=8934,13146,8904,13230,8874,13146 $DEVICE_ID=1001
MM334 202 122 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=12855  $PIN_XY=8934,12852,8904,12855,8874,12852 $DEVICE_ID=1001
MM335 429 202 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=12306  $PIN_XY=8934,12222,8904,12306,8874,12222 $DEVICE_ID=1001
MM336 199 121 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=11931  $PIN_XY=8934,11928,8904,11931,8874,11928 $DEVICE_ID=1001
MM337 GND! 437 212 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=14616  $PIN_XY=8430,14700,8400,14616,8370,14700 $DEVICE_ID=1001
MM338 10 124 437 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=14067  $PIN_XY=8430,14070,8400,14067,8370,14070 $DEVICE_ID=1001
MM339 GND! 433 207 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=13692  $PIN_XY=8430,13776,8400,13692,8370,13776 $DEVICE_ID=1001
MM340 10 123 433 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=13143  $PIN_XY=8430,13146,8400,13143,8370,13146 $DEVICE_ID=1001
MM341 GND! 428 203 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=12768  $PIN_XY=8430,12852,8400,12768,8370,12852 $DEVICE_ID=1001
MM342 10 122 428 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=12219  $PIN_XY=8430,12222,8400,12219,8370,12222 $DEVICE_ID=1001
MM343 GND! 388 200 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=11844  $PIN_XY=8430,11928,8400,11844,8370,11928 $DEVICE_ID=1001
MM344 16 121 391 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=11295  $PIN_XY=10110,11298,10080,11295,10050,11298 $DEVICE_ID=1001
MM345 GND! 398 233 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=10920  $PIN_XY=10110,11004,10080,10920,10050,11004 $DEVICE_ID=1001
MM346 16 120 398 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=10371  $PIN_XY=10110,10374,10080,10371,10050,10374 $DEVICE_ID=1001
MM347 GND! 402 163 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=9996  $PIN_XY=10110,10080,10080,9996,10050,10080 $DEVICE_ID=1001
MM348 16 119 402 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=9447  $PIN_XY=10110,9450,10080,9447,10050,9450 $DEVICE_ID=1001
MM349 GND! 355 162 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=9072  $PIN_XY=10110,9156,10080,9072,10050,9156 $DEVICE_ID=1001
MM350 16 116 355 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=8523  $PIN_XY=10110,8526,10080,8523,10050,8526 $DEVICE_ID=1001
MM351 391 226 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=11382  $PIN_XY=9942,11298,9912,11382,9882,11298 $DEVICE_ID=1001
MM352 233 120 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=11007  $PIN_XY=9942,11004,9912,11007,9882,11004 $DEVICE_ID=1001
MM353 398 233 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=10458  $PIN_XY=9942,10374,9912,10458,9882,10374 $DEVICE_ID=1001
MM354 163 119 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=10083  $PIN_XY=9942,10080,9912,10083,9882,10080 $DEVICE_ID=1001
MM355 402 163 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=9534  $PIN_XY=9942,9450,9912,9534,9882,9450 $DEVICE_ID=1001
MM356 162 116 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=9159  $PIN_XY=9942,9156,9912,9159,9882,9156 $DEVICE_ID=1001
MM357 355 162 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=8610  $PIN_XY=9942,8526,9912,8610,9882,8526 $DEVICE_ID=1001
MM358 8 121 387 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=11295  $PIN_XY=9102,11298,9072,11295,9042,11298 $DEVICE_ID=1001
MM359 GND! 384 197 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=10920  $PIN_XY=9102,11004,9072,10920,9042,11004 $DEVICE_ID=1001
MM360 8 120 384 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=10371  $PIN_XY=9102,10374,9072,10371,9042,10374 $DEVICE_ID=1001
MM361 GND! 382 155 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=9996  $PIN_XY=9102,10080,9072,9996,9042,10080 $DEVICE_ID=1001
MM362 8 119 382 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=9447  $PIN_XY=9102,9450,9072,9447,9042,9450 $DEVICE_ID=1001
MM363 GND! 352 150 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=9072  $PIN_XY=9102,9156,9072,9072,9042,9156 $DEVICE_ID=1001
MM364 8 116 352 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=8523  $PIN_XY=9102,8526,9072,8523,9042,8526 $DEVICE_ID=1001
MM365 387 199 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=11382  $PIN_XY=8934,11298,8904,11382,8874,11298 $DEVICE_ID=1001
MM366 197 120 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=11007  $PIN_XY=8934,11004,8904,11007,8874,11004 $DEVICE_ID=1001
MM367 384 197 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=10458  $PIN_XY=8934,10374,8904,10458,8874,10374 $DEVICE_ID=1001
MM368 155 119 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=10083  $PIN_XY=8934,10080,8904,10083,8874,10080 $DEVICE_ID=1001
MM369 382 155 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=9534  $PIN_XY=8934,9450,8904,9534,8874,9450 $DEVICE_ID=1001
MM370 150 116 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=9159  $PIN_XY=8934,9156,8904,9159,8874,9156 $DEVICE_ID=1001
MM371 352 150 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=8610  $PIN_XY=8934,8526,8904,8610,8874,8526 $DEVICE_ID=1001
MM372 10 121 388 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=11295  $PIN_XY=8430,11298,8400,11295,8370,11298 $DEVICE_ID=1001
MM373 GND! 385 196 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=10920  $PIN_XY=8430,11004,8400,10920,8370,11004 $DEVICE_ID=1001
MM374 10 120 385 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=10371  $PIN_XY=8430,10374,8400,10371,8370,10374 $DEVICE_ID=1001
MM375 GND! 381 154 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=9996  $PIN_XY=8430,10080,8400,9996,8370,10080 $DEVICE_ID=1001
MM376 10 119 381 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=9447  $PIN_XY=8430,9450,8400,9447,8370,9450 $DEVICE_ID=1001
MM377 GND! 351 151 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=9072  $PIN_XY=8430,9156,8400,9072,8370,9156 $DEVICE_ID=1001
MM378 10 116 351 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=8523  $PIN_XY=8430,8526,8400,8523,8370,8526 $DEVICE_ID=1001
MM379 212 124 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=14703  $PIN_XY=8262,14700,8232,14703,8202,14700 $DEVICE_ID=1001
MM380 437 212 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=14154  $PIN_XY=8262,14070,8232,14154,8202,14070 $DEVICE_ID=1001
MM381 207 123 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=13779  $PIN_XY=8262,13776,8232,13779,8202,13776 $DEVICE_ID=1001
MM382 433 207 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=13230  $PIN_XY=8262,13146,8232,13230,8202,13146 $DEVICE_ID=1001
MM383 203 122 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=12855  $PIN_XY=8262,12852,8232,12855,8202,12852 $DEVICE_ID=1001
MM384 428 203 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=12306  $PIN_XY=8262,12222,8232,12306,8202,12222 $DEVICE_ID=1001
MM385 200 121 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=11931  $PIN_XY=8262,11928,8232,11931,8202,11928 $DEVICE_ID=1001
MM386 GND! 438 211 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=14616  $PIN_XY=7758,14700,7728,14616,7698,14700 $DEVICE_ID=1001
MM387 12 124 438 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=14067  $PIN_XY=7758,14070,7728,14067,7698,14070 $DEVICE_ID=1001
MM388 GND! 432 206 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=13692  $PIN_XY=7758,13776,7728,13692,7698,13776 $DEVICE_ID=1001
MM389 12 123 432 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=13143  $PIN_XY=7758,13146,7728,13143,7698,13146 $DEVICE_ID=1001
MM390 GND! 427 204 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=12768  $PIN_XY=7758,12852,7728,12768,7698,12852 $DEVICE_ID=1001
MM391 12 122 427 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=12219  $PIN_XY=7758,12222,7728,12219,7698,12222 $DEVICE_ID=1001
MM392 GND! 389 201 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=11844  $PIN_XY=7758,11928,7728,11844,7698,11928 $DEVICE_ID=1001
MM393 211 124 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=14703  $PIN_XY=7590,14700,7560,14703,7530,14700 $DEVICE_ID=1001
MM394 438 211 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=14154  $PIN_XY=7590,14070,7560,14154,7530,14070 $DEVICE_ID=1001
MM395 206 123 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=13779  $PIN_XY=7590,13776,7560,13779,7530,13776 $DEVICE_ID=1001
MM396 432 206 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=13230  $PIN_XY=7590,13146,7560,13230,7530,13146 $DEVICE_ID=1001
MM397 204 122 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=12855  $PIN_XY=7590,12852,7560,12855,7530,12852 $DEVICE_ID=1001
MM398 427 204 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=12306  $PIN_XY=7590,12222,7560,12306,7530,12222 $DEVICE_ID=1001
MM399 201 121 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=11931  $PIN_XY=7590,11928,7560,11931,7530,11928 $DEVICE_ID=1001
MM400 GND! 435 210 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=14616  $PIN_XY=7086,14700,7056,14616,7026,14700 $DEVICE_ID=1001
MM401 14 124 435 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=14067  $PIN_XY=7086,14070,7056,14067,7026,14070 $DEVICE_ID=1001
MM402 GND! 431 209 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=13692  $PIN_XY=7086,13776,7056,13692,7026,13776 $DEVICE_ID=1001
MM403 14 123 431 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=13143  $PIN_XY=7086,13146,7056,13143,7026,13146 $DEVICE_ID=1001
MM404 GND! 430 205 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=12768  $PIN_XY=7086,12852,7056,12768,7026,12852 $DEVICE_ID=1001
MM405 14 122 430 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=12219  $PIN_XY=7086,12222,7056,12219,7026,12222 $DEVICE_ID=1001
MM406 GND! 390 198 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=11844  $PIN_XY=7086,11928,7056,11844,7026,11928 $DEVICE_ID=1001
MM407 210 124 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=14703  $PIN_XY=6918,14700,6888,14703,6858,14700 $DEVICE_ID=1001
MM408 435 210 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=14154  $PIN_XY=6918,14070,6888,14154,6858,14070 $DEVICE_ID=1001
MM409 209 123 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=13779  $PIN_XY=6918,13776,6888,13779,6858,13776 $DEVICE_ID=1001
MM410 431 209 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=13230  $PIN_XY=6918,13146,6888,13230,6858,13146 $DEVICE_ID=1001
MM411 205 122 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=12855  $PIN_XY=6918,12852,6888,12855,6858,12852 $DEVICE_ID=1001
MM412 430 205 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=12306  $PIN_XY=6918,12222,6888,12306,6858,12222 $DEVICE_ID=1001
MM413 198 121 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=11931  $PIN_XY=6918,11928,6888,11931,6858,11928 $DEVICE_ID=1001
MM414 388 200 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=11382  $PIN_XY=8262,11298,8232,11382,8202,11298 $DEVICE_ID=1001
MM415 196 120 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=11007  $PIN_XY=8262,11004,8232,11007,8202,11004 $DEVICE_ID=1001
MM416 385 196 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=10458  $PIN_XY=8262,10374,8232,10458,8202,10374 $DEVICE_ID=1001
MM417 154 119 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=10083  $PIN_XY=8262,10080,8232,10083,8202,10080 $DEVICE_ID=1001
MM418 381 154 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=9534  $PIN_XY=8262,9450,8232,9534,8202,9450 $DEVICE_ID=1001
MM419 151 116 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=9159  $PIN_XY=8262,9156,8232,9159,8202,9156 $DEVICE_ID=1001
MM420 351 151 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=8610  $PIN_XY=8262,8526,8232,8610,8202,8526 $DEVICE_ID=1001
MM421 12 121 389 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=11295  $PIN_XY=7758,11298,7728,11295,7698,11298 $DEVICE_ID=1001
MM422 GND! 386 195 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=10920  $PIN_XY=7758,11004,7728,10920,7698,11004 $DEVICE_ID=1001
MM423 12 120 386 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=10371  $PIN_XY=7758,10374,7728,10371,7698,10374 $DEVICE_ID=1001
MM424 GND! 380 153 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=9996  $PIN_XY=7758,10080,7728,9996,7698,10080 $DEVICE_ID=1001
MM425 12 119 380 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=9447  $PIN_XY=7758,9450,7728,9447,7698,9450 $DEVICE_ID=1001
MM426 GND! 350 152 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=9072  $PIN_XY=7758,9156,7728,9072,7698,9156 $DEVICE_ID=1001
MM427 12 116 350 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=8523  $PIN_XY=7758,8526,7728,8523,7698,8526 $DEVICE_ID=1001
MM428 389 201 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=11382  $PIN_XY=7590,11298,7560,11382,7530,11298 $DEVICE_ID=1001
MM429 195 120 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=11007  $PIN_XY=7590,11004,7560,11007,7530,11004 $DEVICE_ID=1001
MM430 386 195 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=10458  $PIN_XY=7590,10374,7560,10458,7530,10374 $DEVICE_ID=1001
MM431 153 119 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=10083  $PIN_XY=7590,10080,7560,10083,7530,10080 $DEVICE_ID=1001
MM432 380 153 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=9534  $PIN_XY=7590,9450,7560,9534,7530,9450 $DEVICE_ID=1001
MM433 152 116 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=9159  $PIN_XY=7590,9156,7560,9159,7530,9156 $DEVICE_ID=1001
MM434 350 152 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=8610  $PIN_XY=7590,8526,7560,8610,7530,8526 $DEVICE_ID=1001
MM435 14 121 390 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=11295  $PIN_XY=7086,11298,7056,11295,7026,11298 $DEVICE_ID=1001
MM436 GND! 383 194 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=10920  $PIN_XY=7086,11004,7056,10920,7026,11004 $DEVICE_ID=1001
MM437 14 120 383 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=10371  $PIN_XY=7086,10374,7056,10371,7026,10374 $DEVICE_ID=1001
MM438 GND! 379 157 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=9996  $PIN_XY=7086,10080,7056,9996,7026,10080 $DEVICE_ID=1001
MM439 14 119 379 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=9447  $PIN_XY=7086,9450,7056,9447,7026,9450 $DEVICE_ID=1001
MM440 GND! 354 156 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=9072  $PIN_XY=7086,9156,7056,9072,7026,9156 $DEVICE_ID=1001
MM441 14 116 354 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=8523  $PIN_XY=7086,8526,7056,8523,7026,8526 $DEVICE_ID=1001
MM442 390 198 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=11382  $PIN_XY=6918,11298,6888,11382,6858,11298 $DEVICE_ID=1001
MM443 194 120 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=11007  $PIN_XY=6918,11004,6888,11007,6858,11004 $DEVICE_ID=1001
MM444 383 194 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=10458  $PIN_XY=6918,10374,6888,10458,6858,10374 $DEVICE_ID=1001
MM445 157 119 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=10083  $PIN_XY=6918,10080,6888,10083,6858,10080 $DEVICE_ID=1001
MM446 379 157 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=9534  $PIN_XY=6918,9450,6888,9534,6858,9450 $DEVICE_ID=1001
MM447 156 116 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=9159  $PIN_XY=6918,9156,6888,9159,6858,9156 $DEVICE_ID=1001
MM448 354 156 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=8610  $PIN_XY=6918,8526,6888,8610,6858,8526 $DEVICE_ID=1001
MM449 GND! 371 506 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=8148  $PIN_XY=18174,8232,18144,8148,18114,8232 $DEVICE_ID=1001
MM450 38 115 371 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=7620  $PIN_XY=18174,7602,18144,7620,18114,7602 $DEVICE_ID=1001
MM451 506 115 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=8235  $PIN_XY=18006,8232,17976,8235,17946,8232 $DEVICE_ID=1001
MM452 371 506 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=7707  $PIN_XY=18006,7602,17976,7707,17946,7602 $DEVICE_ID=1001
MM453 GND! 370 505 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=8148  $PIN_XY=17502,8232,17472,8148,17442,8232 $DEVICE_ID=1001
MM454 36 115 370 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=7620  $PIN_XY=17502,7602,17472,7620,17442,7602 $DEVICE_ID=1001
MM455 505 115 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=8235  $PIN_XY=17334,8232,17304,8235,17274,8232 $DEVICE_ID=1001
MM456 370 505 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=7707  $PIN_XY=17334,7602,17304,7707,17274,7602 $DEVICE_ID=1001
MM457 GND! 369 504 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=8148  $PIN_XY=16830,8232,16800,8148,16770,8232 $DEVICE_ID=1001
MM458 34 115 369 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=7620  $PIN_XY=16830,7602,16800,7620,16770,7602 $DEVICE_ID=1001
MM459 504 115 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=8235  $PIN_XY=16662,8232,16632,8235,16602,8232 $DEVICE_ID=1001
MM460 369 504 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=7707  $PIN_XY=16662,7602,16632,7707,16602,7602 $DEVICE_ID=1001
MM461 GND! 368 503 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=8148  $PIN_XY=16158,8232,16128,8148,16098,8232 $DEVICE_ID=1001
MM462 32 115 368 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=7620  $PIN_XY=16158,7602,16128,7620,16098,7602 $DEVICE_ID=1001
MM463 503 115 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=8235  $PIN_XY=15990,8232,15960,8235,15930,8232 $DEVICE_ID=1001
MM464 368 503 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=7707  $PIN_XY=15990,7602,15960,7707,15930,7602 $DEVICE_ID=1001
MM465 GND! 375 507 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=8148  $PIN_XY=15150,8232,15120,8148,15090,8232 $DEVICE_ID=1001
MM466 31 115 375 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=7620  $PIN_XY=15150,7602,15120,7620,15090,7602 $DEVICE_ID=1001
MM467 507 115 30 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=8235  $PIN_XY=14982,8232,14952,8235,14922,8232 $DEVICE_ID=1001
MM468 375 507 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=7707  $PIN_XY=14982,7602,14952,7707,14922,7602 $DEVICE_ID=1001
MM469 GND! 376 508 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=8148  $PIN_XY=14478,8232,14448,8148,14418,8232 $DEVICE_ID=1001
MM470 24 115 376 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=7620  $PIN_XY=14478,7602,14448,7620,14418,7602 $DEVICE_ID=1001
MM471 508 115 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=8235  $PIN_XY=14310,8232,14280,8235,14250,8232 $DEVICE_ID=1001
MM472 376 508 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=7707  $PIN_XY=14310,7602,14280,7707,14250,7602 $DEVICE_ID=1001
MM473 GND! 377 501 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=8148  $PIN_XY=13806,8232,13776,8148,13746,8232 $DEVICE_ID=1001
MM474 26 115 377 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=7620  $PIN_XY=13806,7602,13776,7620,13746,7602 $DEVICE_ID=1001
MM475 501 115 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=8235  $PIN_XY=13638,8232,13608,8235,13578,8232 $DEVICE_ID=1001
MM476 377 501 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=7707  $PIN_XY=13638,7602,13608,7707,13578,7602 $DEVICE_ID=1001
MM477 GND! 378 502 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=8148  $PIN_XY=13134,8232,13104,8148,13074,8232 $DEVICE_ID=1001
MM478 28 115 378 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=7620  $PIN_XY=13134,7602,13104,7620,13074,7602 $DEVICE_ID=1001
MM479 502 115 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=8235  $PIN_XY=12966,8232,12936,8235,12906,8232 $DEVICE_ID=1001
MM480 378 502 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=7707  $PIN_XY=12966,7602,12936,7707,12906,7602 $DEVICE_ID=1001
MM481 GND! 359 497 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=8148  $PIN_XY=12126,8232,12096,8148,12066,8232 $DEVICE_ID=1001
MM482 23 115 359 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=7620  $PIN_XY=12126,7602,12096,7620,12066,7602 $DEVICE_ID=1001
MM483 497 115 22 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=8235  $PIN_XY=11958,8232,11928,8235,11898,8232 $DEVICE_ID=1001
MM484 359 497 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=7707  $PIN_XY=11958,7602,11928,7707,11898,7602 $DEVICE_ID=1001
MM485 GND! 360 498 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=8148  $PIN_XY=11454,8232,11424,8148,11394,8232 $DEVICE_ID=1001
MM486 21 115 360 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=7620  $PIN_XY=11454,7602,11424,7620,11394,7602 $DEVICE_ID=1001
MM487 498 115 20 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=8235  $PIN_XY=11286,8232,11256,8235,11226,8232 $DEVICE_ID=1001
MM488 360 498 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=7707  $PIN_XY=11286,7602,11256,7707,11226,7602 $DEVICE_ID=1001
MM489 GND! 361 499 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=8148  $PIN_XY=10782,8232,10752,8148,10722,8232 $DEVICE_ID=1001
MM490 19 115 361 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=7620  $PIN_XY=10782,7602,10752,7620,10722,7602 $DEVICE_ID=1001
MM491 499 115 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=8235  $PIN_XY=10614,8232,10584,8235,10554,8232 $DEVICE_ID=1001
MM492 361 499 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=7707  $PIN_XY=10614,7602,10584,7707,10554,7602 $DEVICE_ID=1001
MM493 GND! 362 500 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=8148  $PIN_XY=10110,8232,10080,8148,10050,8232 $DEVICE_ID=1001
MM494 16 115 362 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=7620  $PIN_XY=10110,7602,10080,7620,10050,7602 $DEVICE_ID=1001
MM495 500 115 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=8235  $PIN_XY=9942,8232,9912,8235,9882,8232 $DEVICE_ID=1001
MM496 362 500 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=7707  $PIN_XY=9942,7602,9912,7707,9882,7602 $DEVICE_ID=1001
MM497 GND! 347 493 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=8148  $PIN_XY=9102,8232,9072,8148,9042,8232 $DEVICE_ID=1001
MM498 8 115 347 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=7620  $PIN_XY=9102,7602,9072,7620,9042,7602 $DEVICE_ID=1001
MM499 493 115 9 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=8235  $PIN_XY=8934,8232,8904,8235,8874,8232 $DEVICE_ID=1001
MM500 347 493 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=7707  $PIN_XY=8934,7602,8904,7707,8874,7602 $DEVICE_ID=1001
MM501 GND! 348 494 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=8148  $PIN_XY=8430,8232,8400,8148,8370,8232 $DEVICE_ID=1001
MM502 10 115 348 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=7620  $PIN_XY=8430,7602,8400,7620,8370,7602 $DEVICE_ID=1001
MM503 494 115 11 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=8235  $PIN_XY=8262,8232,8232,8235,8202,8232 $DEVICE_ID=1001
MM504 348 494 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=7707  $PIN_XY=8262,7602,8232,7707,8202,7602 $DEVICE_ID=1001
MM505 GND! 349 495 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=8148  $PIN_XY=7758,8232,7728,8148,7698,8232 $DEVICE_ID=1001
MM506 12 115 349 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=7620  $PIN_XY=7758,7602,7728,7620,7698,7602 $DEVICE_ID=1001
MM507 495 115 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=8235  $PIN_XY=7590,8232,7560,8235,7530,8232 $DEVICE_ID=1001
MM508 349 495 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=7707  $PIN_XY=7590,7602,7560,7707,7530,7602 $DEVICE_ID=1001
MM509 GND! 353 496 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=8148  $PIN_XY=7086,8232,7056,8148,7026,8232 $DEVICE_ID=1001
MM510 14 115 353 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=7620  $PIN_XY=7086,7602,7056,7620,7026,7602 $DEVICE_ID=1001
MM511 496 115 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=8235  $PIN_XY=6918,8232,6888,8235,6858,8232 $DEVICE_ID=1001
MM512 353 496 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=7707  $PIN_XY=6918,7602,6888,7707,6858,7602 $DEVICE_ID=1001
MM513 GND! 492 115 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6216 $Y=7686  $PIN_XY=6246,7602,6216,7686,6186,7602 $DEVICE_ID=1001
MM514 115 492 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6048 $Y=7686  $PIN_XY=6078,7602,6048,7686,6018,7602 $DEVICE_ID=1001
MM515 GND! 517 492 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5376 $Y=7707  $PIN_XY=5406,7602,5376,7707,5346,7602 $DEVICE_ID=1001
MM516 492 517 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5208 $Y=7707  $PIN_XY=5238,7602,5208,7707,5178,7602 $DEVICE_ID=1001
MM517 GND! 516 475 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5208 $Y=4935  $PIN_XY=5238,4830,5208,4935,5178,4830 $DEVICE_ID=1001
MM518 475 515 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5040 $Y=4914  $PIN_XY=5070,4830,5040,4914,5010,4830 $DEVICE_ID=1001
MM519 491 514 490 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4704 $Y=7707  $PIN_XY=4734,7602,4704,7707,4674,7602 $DEVICE_ID=1001
MM520 490 A<2> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4536 $Y=7707  $PIN_XY=4566,7602,4536,7707,4506,7602 $DEVICE_ID=1001
MM521 GND! 477 113 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4368 $Y=7203  $PIN_XY=4398,7308,4368,7203,4338,7308 $DEVICE_ID=1001
MM522 GND! 475 114 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4368 $Y=4935  $PIN_XY=4398,4830,4368,4935,4338,4830 $DEVICE_ID=1001
MM523 113 477 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4200 $Y=7203  $PIN_XY=4230,7308,4200,7203,4170,7308 $DEVICE_ID=1001
MM524 114 475 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4200 $Y=4935  $PIN_XY=4230,4830,4200,4935,4170,4830 $DEVICE_ID=1001
MM525 102 478 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3696 $Y=4935  $PIN_XY=3726,4830,3696,4935,3666,4830 $DEVICE_ID=1001
MM526 477 513 476 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=7203  $PIN_XY=3390,7308,3360,7203,3330,7308 $DEVICE_ID=1001
MM527 476 512 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=7203  $PIN_XY=3222,7308,3192,7203,3162,7308 $DEVICE_ID=1001
MM528 478 483 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3192 $Y=4914  $PIN_XY=3222,4830,3192,4914,3162,4830 $DEVICE_ID=1001
MM529 483 484 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2688 $Y=4935  $PIN_XY=2718,4830,2688,4935,2658,4830 $DEVICE_ID=1001
MM530 484 481 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2184 $Y=4935  $PIN_XY=2214,4830,2184,4935,2154,4830 $DEVICE_ID=1001
MM531 481 482 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1680 $Y=4935  $PIN_XY=1710,4830,1680,4935,1650,4830 $DEVICE_ID=1001
MM532 482 479 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1176 $Y=4935  $PIN_XY=1206,4830,1176,4935,1146,4830 $DEVICE_ID=1001
MM533 479 480 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=672 $Y=4935  $PIN_XY=702,4830,672,4935,642,4830 $DEVICE_ID=1001
MM534 480 511 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=168 $Y=4935  $PIN_XY=198,4830,168,4935,138,4830 $DEVICE_ID=1001
MM535 112 144 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17472 $Y=1239  $PIN_XY=17502,1134,17472,1239,17442,1134 $DEVICE_ID=1001
MM536 144 81 489 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16968 $Y=1239  $PIN_XY=16998,1134,16968,1239,16938,1134 $DEVICE_ID=1001
MM537 489 344 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16800 $Y=1218  $PIN_XY=16830,1134,16800,1218,16770,1134 $DEVICE_ID=1001
MM538 GND! 83 344 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=1239  $PIN_XY=16158,1134,16128,1239,16098,1134 $DEVICE_ID=1001
MM539 344 83 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=1239  $PIN_XY=15990,1134,15960,1239,15930,1134 $DEVICE_ID=1001
MM540 111 141 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14448 $Y=1239  $PIN_XY=14478,1134,14448,1239,14418,1134 $DEVICE_ID=1001
MM541 141 85 487 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13944 $Y=1239  $PIN_XY=13974,1134,13944,1239,13914,1134 $DEVICE_ID=1001
MM542 487 345 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13776 $Y=1218  $PIN_XY=13806,1134,13776,1218,13746,1134 $DEVICE_ID=1001
MM543 GND! 87 345 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=1239  $PIN_XY=13134,1134,13104,1239,13074,1134 $DEVICE_ID=1001
MM544 345 87 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=1239  $PIN_XY=12966,1134,12936,1239,12906,1134 $DEVICE_ID=1001
MM545 110 138 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11424 $Y=1239  $PIN_XY=11454,1134,11424,1239,11394,1134 $DEVICE_ID=1001
MM546 138 94 488 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10920 $Y=1239  $PIN_XY=10950,1134,10920,1239,10890,1134 $DEVICE_ID=1001
MM547 488 346 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10752 $Y=1218  $PIN_XY=10782,1134,10752,1218,10722,1134 $DEVICE_ID=1001
MM548 GND! 96 346 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=1239  $PIN_XY=10110,1134,10080,1239,10050,1134 $DEVICE_ID=1001
MM549 346 96 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=1239  $PIN_XY=9942,1134,9912,1239,9882,1134 $DEVICE_ID=1001
MM550 109 135 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8400 $Y=1239  $PIN_XY=8430,1134,8400,1239,8370,1134 $DEVICE_ID=1001
MM551 135 89 486 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7896 $Y=1239  $PIN_XY=7926,1134,7896,1239,7866,1134 $DEVICE_ID=1001
MM552 486 334 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7728 $Y=1218  $PIN_XY=7758,1134,7728,1218,7698,1134 $DEVICE_ID=1001
MM553 GND! 92 334 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=1239  $PIN_XY=7086,1134,7056,1239,7026,1134 $DEVICE_ID=1001
MM554 334 92 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=1239  $PIN_XY=6918,1134,6888,1239,6858,1134 $DEVICE_ID=1001
MM555 107 106 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6384 $Y=1218  $PIN_XY=6414,1134,6384,1218,6354,1134 $DEVICE_ID=1001
MM556 106 WENB 485 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5880 $Y=1218  $PIN_XY=5910,1134,5880,1218,5850,1134 $DEVICE_ID=1001
MM557 485 102 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5712 $Y=1218  $PIN_XY=5742,1134,5712,1218,5682,1134 $DEVICE_ID=1001
MM558 460 273 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=14154  $PIN_XY=18006,14240,17976,14154,17946,14240 $DEVICE_ID=1003
MM559 458 268 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=13230  $PIN_XY=18006,13316,17976,13230,17946,13316 $DEVICE_ID=1003
MM560 453 262 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=12306  $PIN_XY=18006,12392,17976,12306,17946,12392 $DEVICE_ID=1003
MM561 411 259 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=11382  $PIN_XY=18006,11468,17976,11382,17946,11468 $DEVICE_ID=1003
MM562 408 257 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=10458  $PIN_XY=18006,10544,17976,10458,17946,10544 $DEVICE_ID=1003
MM563 406 187 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=9534  $PIN_XY=18006,9620,17976,9534,17946,9620 $DEVICE_ID=1003
MM564 461 272 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=14154  $PIN_XY=17334,14240,17304,14154,17274,14240 $DEVICE_ID=1003
MM565 457 267 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=13230  $PIN_XY=17334,13316,17304,13230,17274,13316 $DEVICE_ID=1003
MM566 452 263 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=12306  $PIN_XY=17334,12392,17304,12306,17274,12392 $DEVICE_ID=1003
MM567 412 260 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=11382  $PIN_XY=17334,11468,17304,11382,17274,11468 $DEVICE_ID=1003
MM568 409 256 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=10458  $PIN_XY=17334,10544,17304,10458,17274,10544 $DEVICE_ID=1003
MM569 405 189 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=9534  $PIN_XY=17334,9620,17304,9534,17274,9620 $DEVICE_ID=1003
MM570 462 271 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=14154  $PIN_XY=16662,14240,16632,14154,16602,14240 $DEVICE_ID=1003
MM571 456 266 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=13230  $PIN_XY=16662,13316,16632,13230,16602,13316 $DEVICE_ID=1003
MM572 451 264 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=12306  $PIN_XY=16662,12392,16632,12306,16602,12392 $DEVICE_ID=1003
MM573 413 261 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=11382  $PIN_XY=16662,11468,16632,11382,16602,11468 $DEVICE_ID=1003
MM574 410 255 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=10458  $PIN_XY=16662,10544,16632,10458,16602,10544 $DEVICE_ID=1003
MM575 404 191 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=9534  $PIN_XY=16662,9620,16632,9534,16602,9620 $DEVICE_ID=1003
MM576 459 270 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=14154  $PIN_XY=15990,14240,15960,14154,15930,14240 $DEVICE_ID=1003
MM577 455 269 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=13230  $PIN_XY=15990,13316,15960,13230,15930,13316 $DEVICE_ID=1003
MM578 454 265 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=12306  $PIN_XY=15990,12392,15960,12306,15930,12392 $DEVICE_ID=1003
MM579 414 258 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=11382  $PIN_XY=15990,11468,15960,11382,15930,11468 $DEVICE_ID=1003
MM580 407 254 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=10458  $PIN_XY=15990,10544,15960,10458,15930,10544 $DEVICE_ID=1003
MM581 403 193 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=9534  $PIN_XY=15990,9620,15960,9534,15930,9620 $DEVICE_ID=1003
MM582 463 234 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=14154  $PIN_XY=14982,14240,14952,14154,14922,14240 $DEVICE_ID=1003
MM583 464 235 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=13230  $PIN_XY=14982,13316,14952,13230,14922,13316 $DEVICE_ID=1003
MM584 465 236 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=12306  $PIN_XY=14982,12392,14952,12306,14922,12392 $DEVICE_ID=1003
MM585 415 237 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=11382  $PIN_XY=14982,11468,14952,11382,14922,11468 $DEVICE_ID=1003
MM586 416 238 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=10458  $PIN_XY=14982,10544,14952,10458,14922,10544 $DEVICE_ID=1003
MM587 417 175 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=9534  $PIN_XY=14982,9620,14952,9534,14922,9620 $DEVICE_ID=1003
MM588 467 240 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=14154  $PIN_XY=14310,14240,14280,14154,14250,14240 $DEVICE_ID=1003
MM589 469 242 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=13230  $PIN_XY=14310,13316,14280,13230,14250,13316 $DEVICE_ID=1003
MM590 473 246 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=12306  $PIN_XY=14310,12392,14280,12306,14250,12392 $DEVICE_ID=1003
MM591 420 250 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=11382  $PIN_XY=14310,11468,14280,11382,14250,11468 $DEVICE_ID=1003
MM592 422 252 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=10458  $PIN_XY=14310,10544,14280,10458,14250,10544 $DEVICE_ID=1003
MM593 424 181 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=9534  $PIN_XY=14310,9620,14280,9534,14250,9620 $DEVICE_ID=1003
MM594 466 239 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=14154  $PIN_XY=13638,14240,13608,14154,13578,14240 $DEVICE_ID=1003
MM595 470 243 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=13230  $PIN_XY=13638,13316,13608,13230,13578,13316 $DEVICE_ID=1003
MM596 474 247 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=12306  $PIN_XY=13638,12392,13608,12306,13578,12392 $DEVICE_ID=1003
MM597 419 249 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=11382  $PIN_XY=13638,11468,13608,11382,13578,11468 $DEVICE_ID=1003
MM598 421 251 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=10458  $PIN_XY=13638,10544,13608,10458,13578,10544 $DEVICE_ID=1003
MM599 425 179 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=9534  $PIN_XY=13638,9620,13608,9534,13578,9620 $DEVICE_ID=1003
MM600 468 241 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=14154  $PIN_XY=12966,14240,12936,14154,12906,14240 $DEVICE_ID=1003
MM601 471 244 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=13230  $PIN_XY=12966,13316,12936,13230,12906,13316 $DEVICE_ID=1003
MM602 472 245 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=12306  $PIN_XY=12966,12392,12936,12306,12906,12392 $DEVICE_ID=1003
MM603 418 248 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=11382  $PIN_XY=12966,11468,12936,11382,12906,11468 $DEVICE_ID=1003
MM604 423 253 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=10458  $PIN_XY=12966,10544,12936,10458,12906,10544 $DEVICE_ID=1003
MM605 426 177 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=9534  $PIN_XY=12966,9620,12936,9534,12906,9620 $DEVICE_ID=1003
MM606 441 216 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=14154  $PIN_XY=11958,14240,11928,14154,11898,14240 $DEVICE_ID=1003
MM607 443 218 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=13230  $PIN_XY=11958,13316,11928,13230,11898,13316 $DEVICE_ID=1003
MM608 448 223 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=12306  $PIN_XY=11958,12392,11928,12306,11898,12392 $DEVICE_ID=1003
MM609 394 229 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=11382  $PIN_XY=11958,11468,11928,11382,11898,11468 $DEVICE_ID=1003
MM610 397 232 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=10458  $PIN_XY=11958,10544,11928,10458,11898,10544 $DEVICE_ID=1003
MM611 399 169 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=9534  $PIN_XY=11958,9620,11928,9534,11898,9620 $DEVICE_ID=1003
MM612 440 215 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=14154  $PIN_XY=11286,14240,11256,14154,11226,14240 $DEVICE_ID=1003
MM613 444 219 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=13230  $PIN_XY=11286,13316,11256,13230,11226,13316 $DEVICE_ID=1003
MM614 449 224 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=12306  $PIN_XY=11286,12392,11256,12306,11226,12392 $DEVICE_ID=1003
MM615 393 228 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=11382  $PIN_XY=11286,11468,11256,11382,11226,11468 $DEVICE_ID=1003
MM616 396 231 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=10458  $PIN_XY=11286,10544,11256,10458,11226,10544 $DEVICE_ID=1003
MM617 400 167 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=9534  $PIN_XY=11286,9620,11256,9534,11226,9620 $DEVICE_ID=1003
MM618 439 214 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=14154  $PIN_XY=10614,14240,10584,14154,10554,14240 $DEVICE_ID=1003
MM619 445 220 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=13230  $PIN_XY=10614,13316,10584,13230,10554,13316 $DEVICE_ID=1003
MM620 450 225 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=12306  $PIN_XY=10614,12392,10584,12306,10554,12392 $DEVICE_ID=1003
MM621 392 227 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=11382  $PIN_XY=10614,11468,10584,11382,10554,11468 $DEVICE_ID=1003
MM622 395 230 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=10458  $PIN_XY=10614,10544,10584,10458,10554,10544 $DEVICE_ID=1003
MM623 401 165 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=9534  $PIN_XY=10614,9620,10584,9534,10554,9620 $DEVICE_ID=1003
MM624 442 217 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=14154  $PIN_XY=9942,14240,9912,14154,9882,14240 $DEVICE_ID=1003
MM625 446 221 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=13230  $PIN_XY=9942,13316,9912,13230,9882,13316 $DEVICE_ID=1003
MM626 447 222 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=12306  $PIN_XY=9942,12392,9912,12306,9882,12392 $DEVICE_ID=1003
MM627 391 226 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=11382  $PIN_XY=9942,11468,9912,11382,9882,11468 $DEVICE_ID=1003
MM628 398 233 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=10458  $PIN_XY=9942,10544,9912,10458,9882,10544 $DEVICE_ID=1003
MM629 402 163 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=9534  $PIN_XY=9942,9620,9912,9534,9882,9620 $DEVICE_ID=1003
MM630 436 213 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=14154  $PIN_XY=8934,14240,8904,14154,8874,14240 $DEVICE_ID=1003
MM631 434 208 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=13230  $PIN_XY=8934,13316,8904,13230,8874,13316 $DEVICE_ID=1003
MM632 429 202 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=12306  $PIN_XY=8934,12392,8904,12306,8874,12392 $DEVICE_ID=1003
MM633 387 199 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=11382  $PIN_XY=8934,11468,8904,11382,8874,11468 $DEVICE_ID=1003
MM634 384 197 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=10458  $PIN_XY=8934,10544,8904,10458,8874,10544 $DEVICE_ID=1003
MM635 382 155 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=9534  $PIN_XY=8934,9620,8904,9534,8874,9620 $DEVICE_ID=1003
MM636 437 212 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=14154  $PIN_XY=8262,14240,8232,14154,8202,14240 $DEVICE_ID=1003
MM637 433 207 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=13230  $PIN_XY=8262,13316,8232,13230,8202,13316 $DEVICE_ID=1003
MM638 428 203 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=12306  $PIN_XY=8262,12392,8232,12306,8202,12392 $DEVICE_ID=1003
MM639 388 200 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=11382  $PIN_XY=8262,11468,8232,11382,8202,11468 $DEVICE_ID=1003
MM640 385 196 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=10458  $PIN_XY=8262,10544,8232,10458,8202,10544 $DEVICE_ID=1003
MM641 381 154 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=9534  $PIN_XY=8262,9620,8232,9534,8202,9620 $DEVICE_ID=1003
MM642 438 211 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=14154  $PIN_XY=7590,14240,7560,14154,7530,14240 $DEVICE_ID=1003
MM643 432 206 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=13230  $PIN_XY=7590,13316,7560,13230,7530,13316 $DEVICE_ID=1003
MM644 427 204 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=12306  $PIN_XY=7590,12392,7560,12306,7530,12392 $DEVICE_ID=1003
MM645 389 201 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=11382  $PIN_XY=7590,11468,7560,11382,7530,11468 $DEVICE_ID=1003
MM646 386 195 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=10458  $PIN_XY=7590,10544,7560,10458,7530,10544 $DEVICE_ID=1003
MM647 380 153 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=9534  $PIN_XY=7590,9620,7560,9534,7530,9620 $DEVICE_ID=1003
MM648 435 210 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=14154  $PIN_XY=6918,14240,6888,14154,6858,14240 $DEVICE_ID=1003
MM649 431 209 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=13230  $PIN_XY=6918,13316,6888,13230,6858,13316 $DEVICE_ID=1003
MM650 430 205 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=12306  $PIN_XY=6918,12392,6888,12306,6858,12392 $DEVICE_ID=1003
MM651 390 198 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=11382  $PIN_XY=6918,11468,6888,11382,6858,11468 $DEVICE_ID=1003
MM652 383 194 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=10458  $PIN_XY=6918,10544,6888,10458,6858,10544 $DEVICE_ID=1003
MM653 379 157 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=9534  $PIN_XY=6918,9620,6888,9534,6858,9620 $DEVICE_ID=1003
MM654 VDD! 75 38 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18312 $Y=7119  $PIN_XY=18342,7138,18312,7119,18282,7138 $DEVICE_ID=1003
MM655 83 185 38 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18312 $Y=6862  $PIN_XY=18342,6848,18312,6862,18282,6848 $DEVICE_ID=1003
MM656 38 75 39 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18144 $Y=7119  $PIN_XY=18174,7138,18144,7119,18114,7138 $DEVICE_ID=1003
MM657 VDD! 97 318 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18144 $Y=3528  $PIN_XY=18174,3442,18144,3528,18114,3442 $DEVICE_ID=1003
MM658 363 186 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=8610  $PIN_XY=18006,8696,17976,8610,17946,8696 $DEVICE_ID=1003
MM659 371 506 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=7707  $PIN_XY=18006,7772,17976,7707,17946,7772 $DEVICE_ID=1003
MM660 39 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=7119  $PIN_XY=18006,7138,17976,7119,17946,7138 $DEVICE_ID=1003
MM661 39 185 81 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17976 $Y=6862  $PIN_XY=18006,6848,17976,6862,17946,6848 $DEVICE_ID=1003
MM662 318 98 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17976 $Y=3549  $PIN_XY=18006,3442,17976,3549,17946,3442 $DEVICE_ID=1003
MM663 VDD! 75 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17640 $Y=7119  $PIN_XY=17670,7138,17640,7119,17610,7138 $DEVICE_ID=1003
MM664 83 184 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17640 $Y=6862  $PIN_XY=17670,6848,17640,6862,17610,6848 $DEVICE_ID=1003
MM665 36 75 37 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17472 $Y=7119  $PIN_XY=17502,7138,17472,7119,17442,7138 $DEVICE_ID=1003
MM666 VDD! 98 317 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=3528  $PIN_XY=17502,3442,17472,3528,17442,3442 $DEVICE_ID=1003
MM667 VDD! 342 82 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=2222  $PIN_XY=17502,2228,17472,2222,17442,2228 $DEVICE_ID=1003
MM668 364 188 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=8610  $PIN_XY=17334,8696,17304,8610,17274,8696 $DEVICE_ID=1003
MM669 370 505 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=7707  $PIN_XY=17334,7772,17304,7707,17274,7772 $DEVICE_ID=1003
MM670 37 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=7119  $PIN_XY=17334,7138,17304,7119,17274,7138 $DEVICE_ID=1003
MM671 37 184 81 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17304 $Y=6862  $PIN_XY=17334,6848,17304,6862,17274,6848 $DEVICE_ID=1003
MM672 317 101 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17304 $Y=3549  $PIN_XY=17334,3442,17304,3549,17274,3442 $DEVICE_ID=1003
MM673 82 342 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17304 $Y=2222  $PIN_XY=17334,2228,17304,2222,17274,2228 $DEVICE_ID=1003
MM674 VDD! 342 82 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17136 $Y=2121  $PIN_XY=17166,2228,17136,2121,17106,2228 $DEVICE_ID=1003
MM675 VDD! 75 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16968 $Y=7119  $PIN_XY=16998,7138,16968,7119,16938,7138 $DEVICE_ID=1003
MM676 83 183 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16968 $Y=6862  $PIN_XY=16998,6848,16968,6862,16938,6848 $DEVICE_ID=1003
MM677 82 342 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16968 $Y=2121  $PIN_XY=16998,2228,16968,2121,16938,2228 $DEVICE_ID=1003
MM678 34 75 35 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16800 $Y=7119  $PIN_XY=16830,7138,16800,7119,16770,7138 $DEVICE_ID=1003
MM679 VDD! 97 316 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16800 $Y=3528  $PIN_XY=16830,3442,16800,3528,16770,3442 $DEVICE_ID=1003
MM680 365 190 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=8610  $PIN_XY=16662,8696,16632,8610,16602,8696 $DEVICE_ID=1003
MM681 369 504 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=7707  $PIN_XY=16662,7772,16632,7707,16602,7772 $DEVICE_ID=1003
MM682 35 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=7119  $PIN_XY=16662,7138,16632,7119,16602,7138 $DEVICE_ID=1003
MM683 35 183 81 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16632 $Y=6862  $PIN_XY=16662,6848,16632,6862,16602,6848 $DEVICE_ID=1003
MM684 316 108 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16632 $Y=3549  $PIN_XY=16662,3442,16632,3549,16602,3442 $DEVICE_ID=1003
MM685 VDD! 343 342 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16632 $Y=2222  $PIN_XY=16662,2228,16632,2222,16602,2228 $DEVICE_ID=1003
MM686 342 343 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16464 $Y=2121  $PIN_XY=16494,2228,16464,2121,16434,2228 $DEVICE_ID=1003
MM687 VDD! 75 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16296 $Y=7119  $PIN_XY=16326,7138,16296,7119,16266,7138 $DEVICE_ID=1003
MM688 83 182 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16296 $Y=6862  $PIN_XY=16326,6848,16296,6862,16266,6848 $DEVICE_ID=1003
MM689 32 75 33 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16128 $Y=7119  $PIN_XY=16158,7138,16128,7119,16098,7138 $DEVICE_ID=1003
MM690 VDD! 108 315 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=3528  $PIN_XY=16158,3442,16128,3528,16098,3442 $DEVICE_ID=1003
MM691 VDD! D<3> 343 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=2222  $PIN_XY=16158,2228,16128,2222,16098,2228 $DEVICE_ID=1003
MM692 366 192 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=8610  $PIN_XY=15990,8696,15960,8610,15930,8696 $DEVICE_ID=1003
MM693 368 503 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=7707  $PIN_XY=15990,7772,15960,7707,15930,7772 $DEVICE_ID=1003
MM694 33 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=7119  $PIN_XY=15990,7138,15960,7119,15930,7138 $DEVICE_ID=1003
MM695 33 182 81 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15960 $Y=6862  $PIN_XY=15990,6848,15960,6862,15930,6848 $DEVICE_ID=1003
MM696 315 101 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=3549  $PIN_XY=15990,3442,15960,3549,15930,3442 $DEVICE_ID=1003
MM697 343 D<3> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=2121  $PIN_XY=15990,2228,15960,2121,15930,2228 $DEVICE_ID=1003
MM698 VDD! 75 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15288 $Y=7119  $PIN_XY=15318,7138,15288,7119,15258,7138 $DEVICE_ID=1003
MM699 87 170 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15288 $Y=6862  $PIN_XY=15318,6848,15288,6862,15258,6848 $DEVICE_ID=1003
MM700 31 75 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=15120 $Y=7119  $PIN_XY=15150,7138,15120,7119,15090,7138 $DEVICE_ID=1003
MM701 VDD! 97 322 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15120 $Y=3528  $PIN_XY=15150,3442,15120,3528,15090,3442 $DEVICE_ID=1003
MM702 367 174 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=8610  $PIN_XY=14982,8696,14952,8610,14922,8696 $DEVICE_ID=1003
MM703 375 507 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=7707  $PIN_XY=14982,7772,14952,7707,14922,7772 $DEVICE_ID=1003
MM704 30 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=7119  $PIN_XY=14982,7138,14952,7119,14922,7138 $DEVICE_ID=1003
MM705 30 170 85 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14952 $Y=6862  $PIN_XY=14982,6848,14952,6862,14922,6848 $DEVICE_ID=1003
MM706 322 98 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14952 $Y=3549  $PIN_XY=14982,3442,14952,3549,14922,3442 $DEVICE_ID=1003
MM707 VDD! 75 24 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14616 $Y=7119  $PIN_XY=14646,7138,14616,7119,14586,7138 $DEVICE_ID=1003
MM708 87 171 24 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14616 $Y=6862  $PIN_XY=14646,6848,14616,6862,14586,6848 $DEVICE_ID=1003
MM709 24 75 25 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14448 $Y=7119  $PIN_XY=14478,7138,14448,7119,14418,7138 $DEVICE_ID=1003
MM710 VDD! 98 321 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=3528  $PIN_XY=14478,3442,14448,3528,14418,3442 $DEVICE_ID=1003
MM711 VDD! 339 86 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=2222  $PIN_XY=14478,2228,14448,2222,14418,2228 $DEVICE_ID=1003
MM712 374 180 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=8610  $PIN_XY=14310,8696,14280,8610,14250,8696 $DEVICE_ID=1003
MM713 376 508 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=7707  $PIN_XY=14310,7772,14280,7707,14250,7772 $DEVICE_ID=1003
MM714 25 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=7119  $PIN_XY=14310,7138,14280,7119,14250,7138 $DEVICE_ID=1003
MM715 25 171 85 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14280 $Y=6862  $PIN_XY=14310,6848,14280,6862,14250,6848 $DEVICE_ID=1003
MM716 321 101 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14280 $Y=3549  $PIN_XY=14310,3442,14280,3549,14250,3442 $DEVICE_ID=1003
MM717 86 339 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14280 $Y=2222  $PIN_XY=14310,2228,14280,2222,14250,2228 $DEVICE_ID=1003
MM718 VDD! 339 86 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14112 $Y=2121  $PIN_XY=14142,2228,14112,2121,14082,2228 $DEVICE_ID=1003
MM719 VDD! 75 26 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13944 $Y=7119  $PIN_XY=13974,7138,13944,7119,13914,7138 $DEVICE_ID=1003
MM720 87 172 26 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13944 $Y=6862  $PIN_XY=13974,6848,13944,6862,13914,6848 $DEVICE_ID=1003
MM721 86 339 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13944 $Y=2121  $PIN_XY=13974,2228,13944,2121,13914,2228 $DEVICE_ID=1003
MM722 26 75 27 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13776 $Y=7119  $PIN_XY=13806,7138,13776,7119,13746,7138 $DEVICE_ID=1003
MM723 VDD! 97 320 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13776 $Y=3528  $PIN_XY=13806,3442,13776,3528,13746,3442 $DEVICE_ID=1003
MM724 373 178 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=8610  $PIN_XY=13638,8696,13608,8610,13578,8696 $DEVICE_ID=1003
MM725 377 501 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=7707  $PIN_XY=13638,7772,13608,7707,13578,7772 $DEVICE_ID=1003
MM726 27 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=7119  $PIN_XY=13638,7138,13608,7119,13578,7138 $DEVICE_ID=1003
MM727 27 172 85 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13608 $Y=6862  $PIN_XY=13638,6848,13608,6862,13578,6848 $DEVICE_ID=1003
MM728 320 108 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13608 $Y=3549  $PIN_XY=13638,3442,13608,3549,13578,3442 $DEVICE_ID=1003
MM729 VDD! 340 339 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13608 $Y=2222  $PIN_XY=13638,2228,13608,2222,13578,2228 $DEVICE_ID=1003
MM730 339 340 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13440 $Y=2121  $PIN_XY=13470,2228,13440,2121,13410,2228 $DEVICE_ID=1003
MM731 VDD! 75 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13272 $Y=7119  $PIN_XY=13302,7138,13272,7119,13242,7138 $DEVICE_ID=1003
MM732 87 173 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13272 $Y=6862  $PIN_XY=13302,6848,13272,6862,13242,6848 $DEVICE_ID=1003
MM733 28 75 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13104 $Y=7119  $PIN_XY=13134,7138,13104,7119,13074,7138 $DEVICE_ID=1003
MM734 VDD! 108 319 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=3528  $PIN_XY=13134,3442,13104,3528,13074,3442 $DEVICE_ID=1003
MM735 VDD! D<2> 340 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=2222  $PIN_XY=13134,2228,13104,2222,13074,2228 $DEVICE_ID=1003
MM736 372 176 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=8610  $PIN_XY=12966,8696,12936,8610,12906,8696 $DEVICE_ID=1003
MM737 378 502 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=7707  $PIN_XY=12966,7772,12936,7707,12906,7772 $DEVICE_ID=1003
MM738 29 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=7119  $PIN_XY=12966,7138,12936,7119,12906,7138 $DEVICE_ID=1003
MM739 29 173 85 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12936 $Y=6862  $PIN_XY=12966,6848,12936,6862,12906,6848 $DEVICE_ID=1003
MM740 319 101 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=3549  $PIN_XY=12966,3442,12936,3549,12906,3442 $DEVICE_ID=1003
MM741 340 D<2> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=2121  $PIN_XY=12966,2228,12936,2121,12906,2228 $DEVICE_ID=1003
MM742 VDD! 75 23 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12264 $Y=7119  $PIN_XY=12294,7138,12264,7119,12234,7138 $DEVICE_ID=1003
MM743 96 158 23 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12264 $Y=6862  $PIN_XY=12294,6848,12264,6862,12234,6848 $DEVICE_ID=1003
MM744 23 75 22 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=12096 $Y=7119  $PIN_XY=12126,7138,12096,7119,12066,7138 $DEVICE_ID=1003
MM745 VDD! 97 330 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12096 $Y=3528  $PIN_XY=12126,3442,12096,3528,12066,3442 $DEVICE_ID=1003
MM746 358 168 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=8610  $PIN_XY=11958,8696,11928,8610,11898,8696 $DEVICE_ID=1003
MM747 359 497 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=7707  $PIN_XY=11958,7772,11928,7707,11898,7772 $DEVICE_ID=1003
MM748 22 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=7119  $PIN_XY=11958,7138,11928,7119,11898,7138 $DEVICE_ID=1003
MM749 22 158 94 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11928 $Y=6862  $PIN_XY=11958,6848,11928,6862,11898,6848 $DEVICE_ID=1003
MM750 330 98 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11928 $Y=3549  $PIN_XY=11958,3442,11928,3549,11898,3442 $DEVICE_ID=1003
MM751 VDD! 75 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11592 $Y=7119  $PIN_XY=11622,7138,11592,7119,11562,7138 $DEVICE_ID=1003
MM752 96 159 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11592 $Y=6862  $PIN_XY=11622,6848,11592,6862,11562,6848 $DEVICE_ID=1003
MM753 21 75 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11424 $Y=7119  $PIN_XY=11454,7138,11424,7119,11394,7138 $DEVICE_ID=1003
MM754 VDD! 98 329 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=3528  $PIN_XY=11454,3442,11424,3528,11394,3442 $DEVICE_ID=1003
MM755 VDD! 336 95 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=2222  $PIN_XY=11454,2228,11424,2222,11394,2228 $DEVICE_ID=1003
MM756 357 166 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=8610  $PIN_XY=11286,8696,11256,8610,11226,8696 $DEVICE_ID=1003
MM757 360 498 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=7707  $PIN_XY=11286,7772,11256,7707,11226,7772 $DEVICE_ID=1003
MM758 20 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=7119  $PIN_XY=11286,7138,11256,7119,11226,7138 $DEVICE_ID=1003
MM759 20 159 94 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11256 $Y=6862  $PIN_XY=11286,6848,11256,6862,11226,6848 $DEVICE_ID=1003
MM760 329 101 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11256 $Y=3549  $PIN_XY=11286,3442,11256,3549,11226,3442 $DEVICE_ID=1003
MM761 95 336 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11256 $Y=2222  $PIN_XY=11286,2228,11256,2222,11226,2228 $DEVICE_ID=1003
MM762 VDD! 336 95 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11088 $Y=2121  $PIN_XY=11118,2228,11088,2121,11058,2228 $DEVICE_ID=1003
MM763 VDD! 75 19 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10920 $Y=7119  $PIN_XY=10950,7138,10920,7119,10890,7138 $DEVICE_ID=1003
MM764 96 160 19 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10920 $Y=6862  $PIN_XY=10950,6848,10920,6862,10890,6848 $DEVICE_ID=1003
MM765 95 336 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10920 $Y=2121  $PIN_XY=10950,2228,10920,2121,10890,2228 $DEVICE_ID=1003
MM766 19 75 18 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10752 $Y=7119  $PIN_XY=10782,7138,10752,7119,10722,7138 $DEVICE_ID=1003
MM767 VDD! 97 328 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10752 $Y=3528  $PIN_XY=10782,3442,10752,3528,10722,3442 $DEVICE_ID=1003
MM768 356 164 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=8610  $PIN_XY=10614,8696,10584,8610,10554,8696 $DEVICE_ID=1003
MM769 361 499 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=7707  $PIN_XY=10614,7772,10584,7707,10554,7772 $DEVICE_ID=1003
MM770 18 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=7119  $PIN_XY=10614,7138,10584,7119,10554,7138 $DEVICE_ID=1003
MM771 18 160 94 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10584 $Y=6862  $PIN_XY=10614,6848,10584,6862,10554,6848 $DEVICE_ID=1003
MM772 328 108 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10584 $Y=3549  $PIN_XY=10614,3442,10584,3549,10554,3442 $DEVICE_ID=1003
MM773 VDD! 337 336 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10584 $Y=2222  $PIN_XY=10614,2228,10584,2222,10554,2228 $DEVICE_ID=1003
MM774 336 337 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10416 $Y=2121  $PIN_XY=10446,2228,10416,2121,10386,2228 $DEVICE_ID=1003
MM775 VDD! 75 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10248 $Y=7119  $PIN_XY=10278,7138,10248,7119,10218,7138 $DEVICE_ID=1003
MM776 96 161 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10248 $Y=6862  $PIN_XY=10278,6848,10248,6862,10218,6848 $DEVICE_ID=1003
MM777 16 75 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10080 $Y=7119  $PIN_XY=10110,7138,10080,7119,10050,7138 $DEVICE_ID=1003
MM778 VDD! 108 327 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=3528  $PIN_XY=10110,3442,10080,3528,10050,3442 $DEVICE_ID=1003
MM779 VDD! D<1> 337 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=2222  $PIN_XY=10110,2228,10080,2222,10050,2228 $DEVICE_ID=1003
MM780 355 162 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=8610  $PIN_XY=9942,8696,9912,8610,9882,8696 $DEVICE_ID=1003
MM781 362 500 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=7707  $PIN_XY=9942,7772,9912,7707,9882,7772 $DEVICE_ID=1003
MM782 17 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=7119  $PIN_XY=9942,7138,9912,7119,9882,7138 $DEVICE_ID=1003
MM783 17 161 94 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9912 $Y=6862  $PIN_XY=9942,6848,9912,6862,9882,6848 $DEVICE_ID=1003
MM784 327 101 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=3549  $PIN_XY=9942,3442,9912,3549,9882,3442 $DEVICE_ID=1003
MM785 337 D<1> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=2121  $PIN_XY=9942,2228,9912,2121,9882,2228 $DEVICE_ID=1003
MM786 VDD! 75 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9240 $Y=7119  $PIN_XY=9270,7138,9240,7119,9210,7138 $DEVICE_ID=1003
MM787 92 146 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9240 $Y=6862  $PIN_XY=9270,6848,9240,6862,9210,6848 $DEVICE_ID=1003
MM788 8 75 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9072 $Y=7119  $PIN_XY=9102,7138,9072,7119,9042,7138 $DEVICE_ID=1003
MM789 VDD! 97 326 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9072 $Y=3528  $PIN_XY=9102,3442,9072,3528,9042,3442 $DEVICE_ID=1003
MM790 352 150 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=8610  $PIN_XY=8934,8696,8904,8610,8874,8696 $DEVICE_ID=1003
MM791 347 493 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=7707  $PIN_XY=8934,7772,8904,7707,8874,7772 $DEVICE_ID=1003
MM792 9 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=7119  $PIN_XY=8934,7138,8904,7119,8874,7138 $DEVICE_ID=1003
MM793 9 146 89 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8904 $Y=6862  $PIN_XY=8934,6848,8904,6862,8874,6848 $DEVICE_ID=1003
MM794 326 98 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8904 $Y=3549  $PIN_XY=8934,3442,8904,3549,8874,3442 $DEVICE_ID=1003
MM795 VDD! 75 10 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8568 $Y=7119  $PIN_XY=8598,7138,8568,7119,8538,7138 $DEVICE_ID=1003
MM796 92 147 10 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8568 $Y=6862  $PIN_XY=8598,6848,8568,6862,8538,6848 $DEVICE_ID=1003
MM797 10 75 11 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8400 $Y=7119  $PIN_XY=8430,7138,8400,7119,8370,7138 $DEVICE_ID=1003
MM798 VDD! 98 325 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=3528  $PIN_XY=8430,3442,8400,3528,8370,3442 $DEVICE_ID=1003
MM799 VDD! 332 91 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=2222  $PIN_XY=8430,2228,8400,2222,8370,2228 $DEVICE_ID=1003
MM800 351 151 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=8610  $PIN_XY=8262,8696,8232,8610,8202,8696 $DEVICE_ID=1003
MM801 348 494 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=7707  $PIN_XY=8262,7772,8232,7707,8202,7772 $DEVICE_ID=1003
MM802 11 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=7119  $PIN_XY=8262,7138,8232,7119,8202,7138 $DEVICE_ID=1003
MM803 11 147 89 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8232 $Y=6862  $PIN_XY=8262,6848,8232,6862,8202,6848 $DEVICE_ID=1003
MM804 325 101 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8232 $Y=3549  $PIN_XY=8262,3442,8232,3549,8202,3442 $DEVICE_ID=1003
MM805 91 332 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8232 $Y=2222  $PIN_XY=8262,2228,8232,2222,8202,2228 $DEVICE_ID=1003
MM806 VDD! 332 91 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8064 $Y=2121  $PIN_XY=8094,2228,8064,2121,8034,2228 $DEVICE_ID=1003
MM807 VDD! 75 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7896 $Y=7119  $PIN_XY=7926,7138,7896,7119,7866,7138 $DEVICE_ID=1003
MM808 92 148 12 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7896 $Y=6862  $PIN_XY=7926,6848,7896,6862,7866,6848 $DEVICE_ID=1003
MM809 91 332 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7896 $Y=2121  $PIN_XY=7926,2228,7896,2121,7866,2228 $DEVICE_ID=1003
MM810 12 75 13 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7728 $Y=7119  $PIN_XY=7758,7138,7728,7119,7698,7138 $DEVICE_ID=1003
MM811 VDD! 97 324 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7728 $Y=3528  $PIN_XY=7758,3442,7728,3528,7698,3442 $DEVICE_ID=1003
MM812 350 152 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=8610  $PIN_XY=7590,8696,7560,8610,7530,8696 $DEVICE_ID=1003
MM813 349 495 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=7707  $PIN_XY=7590,7772,7560,7707,7530,7772 $DEVICE_ID=1003
MM814 13 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=7119  $PIN_XY=7590,7138,7560,7119,7530,7138 $DEVICE_ID=1003
MM815 13 148 89 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7560 $Y=6862  $PIN_XY=7590,6848,7560,6862,7530,6848 $DEVICE_ID=1003
MM816 324 108 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7560 $Y=3549  $PIN_XY=7590,3442,7560,3549,7530,3442 $DEVICE_ID=1003
MM817 VDD! 333 332 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7560 $Y=2222  $PIN_XY=7590,2228,7560,2222,7530,2228 $DEVICE_ID=1003
MM818 332 333 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7392 $Y=2121  $PIN_XY=7422,2228,7392,2121,7362,2228 $DEVICE_ID=1003
MM819 VDD! 75 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7224 $Y=7119  $PIN_XY=7254,7138,7224,7119,7194,7138 $DEVICE_ID=1003
MM820 92 149 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7224 $Y=6862  $PIN_XY=7254,6848,7224,6862,7194,6848 $DEVICE_ID=1003
MM821 14 75 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7056 $Y=7119  $PIN_XY=7086,7138,7056,7119,7026,7138 $DEVICE_ID=1003
MM822 VDD! 108 323 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=3528  $PIN_XY=7086,3442,7056,3528,7026,3442 $DEVICE_ID=1003
MM823 VDD! D<0> 333 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=2222  $PIN_XY=7086,2228,7056,2222,7026,2228 $DEVICE_ID=1003
MM824 354 156 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=8610  $PIN_XY=6918,8696,6888,8610,6858,8696 $DEVICE_ID=1003
MM825 353 496 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=7707  $PIN_XY=6918,7772,6888,7707,6858,7772 $DEVICE_ID=1003
MM826 15 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=7119  $PIN_XY=6918,7138,6888,7119,6858,7138 $DEVICE_ID=1003
MM827 15 149 89 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6888 $Y=6862  $PIN_XY=6918,6848,6888,6862,6858,6848 $DEVICE_ID=1003
MM828 323 101 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=3549  $PIN_XY=6918,3442,6888,3549,6858,3442 $DEVICE_ID=1003
MM829 333 D<0> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=2121  $PIN_XY=6918,2228,6888,2121,6858,2228 $DEVICE_ID=1003
MM830 VDD! 313 117 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6552 $Y=6842  $PIN_XY=6582,6848,6552,6842,6522,6848 $DEVICE_ID=1003
MM831 VDD! 314 101 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6552 $Y=3528  $PIN_XY=6582,3442,6552,3528,6522,3442 $DEVICE_ID=1003
MM832 117 313 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6384 $Y=6762  $PIN_XY=6414,6848,6384,6762,6354,6848 $DEVICE_ID=1003
MM833 101 314 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6384 $Y=3448  $PIN_XY=6414,3442,6384,3448,6354,3442 $DEVICE_ID=1003
MM834 VDD! 113 314 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6048 $Y=3528  $PIN_XY=6078,3442,6048,3528,6018,3442 $DEVICE_ID=1003
MM835 313 103 312 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5880 $Y=6741  $PIN_XY=5910,6848,5880,6741,5850,6848 $DEVICE_ID=1003
MM836 314 WS0BAR VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5880 $Y=3549  $PIN_XY=5910,3442,5880,3549,5850,3442 $DEVICE_ID=1003
MM837 312 114 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5712 $Y=6762  $PIN_XY=5742,6848,5712,6762,5682,6848 $DEVICE_ID=1003
MM838 VDD! 308 WS0BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5376 $Y=4070  $PIN_XY=5406,4076,5376,4070,5346,4076 $DEVICE_ID=1003
MM839 WS0BAR 308 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5208 $Y=4070  $PIN_XY=5238,4076,5208,4070,5178,4076 $DEVICE_ID=1003
MM840 VDD! 308 WS0BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5040 $Y=3969  $PIN_XY=5070,4076,5040,3969,5010,4076 $DEVICE_ID=1003
MM841 WS0BAR 308 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4872 $Y=3969  $PIN_XY=4902,4076,4872,3969,4842,4076 $DEVICE_ID=1003
MM842 VDD! 509 308 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4368 $Y=3969  $PIN_XY=4398,4076,4368,3969,4338,4076 $DEVICE_ID=1003
MM843 308 305 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4200 $Y=3969  $PIN_XY=4230,4076,4200,3969,4170,4076 $DEVICE_ID=1003
MM844 VDD! 310 305 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3360 $Y=4070  $PIN_XY=3390,4076,3360,4070,3330,4076 $DEVICE_ID=1003
MM845 305 310 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3192 $Y=3990  $PIN_XY=3222,4076,3192,3990,3162,4076 $DEVICE_ID=1003
MM846 VDD! 311 310 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2856 $Y=4070  $PIN_XY=2886,4076,2856,4070,2826,4076 $DEVICE_ID=1003
MM847 310 311 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2688 $Y=3969  $PIN_XY=2718,4076,2688,3969,2658,4076 $DEVICE_ID=1003
MM848 VDD! 309 311 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2184 $Y=3969  $PIN_XY=2214,4076,2184,3969,2154,4076 $DEVICE_ID=1003
MM849 311 A<0> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2016 $Y=3969  $PIN_XY=2046,4076,2016,3969,1986,4076 $DEVICE_ID=1003
MM850 VDD! WENB 309 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1680 $Y=4070  $PIN_XY=1710,4076,1680,4070,1650,4076 $DEVICE_ID=1003
MM851 309 WENB VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1512 $Y=3990  $PIN_XY=1542,4076,1512,3990,1482,4076 $DEVICE_ID=1003
MM852 VDD! 341 80 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=18312 $Y=1600  $PIN_XY=18342,1594,18312,1600,18282,1594 $DEVICE_ID=1003
MM853 80 341 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18144 $Y=1600  $PIN_XY=18174,1594,18144,1600,18114,1594 $DEVICE_ID=1003
MM854 VDD! 341 80 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17976 $Y=1680  $PIN_XY=18006,1594,17976,1680,17946,1594 $DEVICE_ID=1003
MM855 80 341 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17808 $Y=1680  $PIN_XY=17838,1594,17808,1680,17778,1594 $DEVICE_ID=1003
MM856 VDD! 144 112 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17640 $Y=1298  $PIN_XY=17670,1304,17640,1298,17610,1304 $DEVICE_ID=1003
MM857 VDD! 145 341 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=17472 $Y=1579  $PIN_XY=17502,1594,17472,1579,17442,1594 $DEVICE_ID=1003
MM858 112 144 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=17472 $Y=1239  $PIN_XY=17502,1304,17472,1239,17442,1304 $DEVICE_ID=1003
MM859 341 145 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17304 $Y=1600  $PIN_XY=17334,1594,17304,1600,17274,1594 $DEVICE_ID=1003
MM860 VDD! 145 341 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17136 $Y=1701  $PIN_XY=17166,1594,17136,1701,17106,1594 $DEVICE_ID=1003
MM861 341 145 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16968 $Y=1680  $PIN_XY=16998,1594,16968,1680,16938,1594 $DEVICE_ID=1003
MM862 VDD! 81 144 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16968 $Y=1239  $PIN_XY=16998,1304,16968,1239,16938,1304 $DEVICE_ID=1003
MM863 144 344 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16800 $Y=1218  $PIN_XY=16830,1304,16800,1218,16770,1304 $DEVICE_ID=1003
MM864 VDD! 143 145 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16632 $Y=1600  $PIN_XY=16662,1594,16632,1600,16602,1594 $DEVICE_ID=1003
MM865 145 143 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=16464 $Y=1680  $PIN_XY=16494,1594,16464,1680,16434,1594 $DEVICE_ID=1003
MM866 VDD! 83 344 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16464 $Y=1319  $PIN_XY=16494,1304,16464,1319,16434,1304 $DEVICE_ID=1003
MM867 344 83 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16296 $Y=1298  $PIN_XY=16326,1304,16296,1298,16266,1304 $DEVICE_ID=1003
MM868 VDD! D<3> 143 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=16128 $Y=1579  $PIN_XY=16158,1594,16128,1579,16098,1594 $DEVICE_ID=1003
MM869 VDD! 83 344 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16128 $Y=1239  $PIN_XY=16158,1304,16128,1239,16098,1304 $DEVICE_ID=1003
MM870 143 D<3> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=1680  $PIN_XY=15990,1594,15960,1680,15930,1594 $DEVICE_ID=1003
MM871 344 83 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=15960 $Y=1239  $PIN_XY=15990,1304,15960,1239,15930,1304 $DEVICE_ID=1003
MM872 VDD! 338 84 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=15288 $Y=1600  $PIN_XY=15318,1594,15288,1600,15258,1594 $DEVICE_ID=1003
MM873 84 338 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=15120 $Y=1600  $PIN_XY=15150,1594,15120,1600,15090,1594 $DEVICE_ID=1003
MM874 VDD! 338 84 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14952 $Y=1680  $PIN_XY=14982,1594,14952,1680,14922,1594 $DEVICE_ID=1003
MM875 84 338 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14784 $Y=1680  $PIN_XY=14814,1594,14784,1680,14754,1594 $DEVICE_ID=1003
MM876 VDD! 141 111 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14616 $Y=1298  $PIN_XY=14646,1304,14616,1298,14586,1304 $DEVICE_ID=1003
MM877 VDD! 142 338 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=14448 $Y=1579  $PIN_XY=14478,1594,14448,1579,14418,1594 $DEVICE_ID=1003
MM878 111 141 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=14448 $Y=1239  $PIN_XY=14478,1304,14448,1239,14418,1304 $DEVICE_ID=1003
MM879 338 142 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14280 $Y=1600  $PIN_XY=14310,1594,14280,1600,14250,1594 $DEVICE_ID=1003
MM880 VDD! 142 338 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14112 $Y=1701  $PIN_XY=14142,1594,14112,1701,14082,1594 $DEVICE_ID=1003
MM881 338 142 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13944 $Y=1680  $PIN_XY=13974,1594,13944,1680,13914,1594 $DEVICE_ID=1003
MM882 VDD! 85 141 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13944 $Y=1239  $PIN_XY=13974,1304,13944,1239,13914,1304 $DEVICE_ID=1003
MM883 141 345 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13776 $Y=1218  $PIN_XY=13806,1304,13776,1218,13746,1304 $DEVICE_ID=1003
MM884 VDD! 140 142 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13608 $Y=1600  $PIN_XY=13638,1594,13608,1600,13578,1594 $DEVICE_ID=1003
MM885 142 140 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=13440 $Y=1680  $PIN_XY=13470,1594,13440,1680,13410,1594 $DEVICE_ID=1003
MM886 VDD! 87 345 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13440 $Y=1319  $PIN_XY=13470,1304,13440,1319,13410,1304 $DEVICE_ID=1003
MM887 345 87 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13272 $Y=1298  $PIN_XY=13302,1304,13272,1298,13242,1304 $DEVICE_ID=1003
MM888 VDD! D<2> 140 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=13104 $Y=1579  $PIN_XY=13134,1594,13104,1579,13074,1594 $DEVICE_ID=1003
MM889 VDD! 87 345 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13104 $Y=1239  $PIN_XY=13134,1304,13104,1239,13074,1304 $DEVICE_ID=1003
MM890 140 D<2> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=1680  $PIN_XY=12966,1594,12936,1680,12906,1594 $DEVICE_ID=1003
MM891 345 87 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=12936 $Y=1239  $PIN_XY=12966,1304,12936,1239,12906,1304 $DEVICE_ID=1003
MM892 VDD! 335 93 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=12264 $Y=1600  $PIN_XY=12294,1594,12264,1600,12234,1594 $DEVICE_ID=1003
MM893 93 335 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=12096 $Y=1600  $PIN_XY=12126,1594,12096,1600,12066,1594 $DEVICE_ID=1003
MM894 VDD! 335 93 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11928 $Y=1680  $PIN_XY=11958,1594,11928,1680,11898,1594 $DEVICE_ID=1003
MM895 93 335 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11760 $Y=1680  $PIN_XY=11790,1594,11760,1680,11730,1594 $DEVICE_ID=1003
MM896 VDD! 138 110 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11592 $Y=1298  $PIN_XY=11622,1304,11592,1298,11562,1304 $DEVICE_ID=1003
MM897 VDD! 139 335 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=11424 $Y=1579  $PIN_XY=11454,1594,11424,1579,11394,1594 $DEVICE_ID=1003
MM898 110 138 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=11424 $Y=1239  $PIN_XY=11454,1304,11424,1239,11394,1304 $DEVICE_ID=1003
MM899 335 139 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11256 $Y=1600  $PIN_XY=11286,1594,11256,1600,11226,1594 $DEVICE_ID=1003
MM900 VDD! 139 335 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11088 $Y=1701  $PIN_XY=11118,1594,11088,1701,11058,1594 $DEVICE_ID=1003
MM901 335 139 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10920 $Y=1680  $PIN_XY=10950,1594,10920,1680,10890,1594 $DEVICE_ID=1003
MM902 VDD! 94 138 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10920 $Y=1239  $PIN_XY=10950,1304,10920,1239,10890,1304 $DEVICE_ID=1003
MM903 138 346 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10752 $Y=1218  $PIN_XY=10782,1304,10752,1218,10722,1304 $DEVICE_ID=1003
MM904 VDD! 137 139 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10584 $Y=1600  $PIN_XY=10614,1594,10584,1600,10554,1594 $DEVICE_ID=1003
MM905 139 137 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=10416 $Y=1680  $PIN_XY=10446,1594,10416,1680,10386,1594 $DEVICE_ID=1003
MM906 VDD! 96 346 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10416 $Y=1319  $PIN_XY=10446,1304,10416,1319,10386,1304 $DEVICE_ID=1003
MM907 346 96 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10248 $Y=1298  $PIN_XY=10278,1304,10248,1298,10218,1304 $DEVICE_ID=1003
MM908 VDD! D<1> 137 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=10080 $Y=1579  $PIN_XY=10110,1594,10080,1579,10050,1594 $DEVICE_ID=1003
MM909 VDD! 96 346 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10080 $Y=1239  $PIN_XY=10110,1304,10080,1239,10050,1304 $DEVICE_ID=1003
MM910 137 D<1> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=1680  $PIN_XY=9942,1594,9912,1680,9882,1594 $DEVICE_ID=1003
MM911 346 96 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=9912 $Y=1239  $PIN_XY=9942,1304,9912,1239,9882,1304 $DEVICE_ID=1003
MM912 VDD! 331 88 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9240 $Y=1600  $PIN_XY=9270,1594,9240,1600,9210,1594 $DEVICE_ID=1003
MM913 88 331 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9072 $Y=1600  $PIN_XY=9102,1594,9072,1600,9042,1594 $DEVICE_ID=1003
MM914 VDD! 331 88 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8904 $Y=1680  $PIN_XY=8934,1594,8904,1680,8874,1594 $DEVICE_ID=1003
MM915 88 331 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8736 $Y=1680  $PIN_XY=8766,1594,8736,1680,8706,1594 $DEVICE_ID=1003
MM916 VDD! 135 109 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8568 $Y=1298  $PIN_XY=8598,1304,8568,1298,8538,1304 $DEVICE_ID=1003
MM917 VDD! 136 331 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8400 $Y=1579  $PIN_XY=8430,1594,8400,1579,8370,1594 $DEVICE_ID=1003
MM918 109 135 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8400 $Y=1239  $PIN_XY=8430,1304,8400,1239,8370,1304 $DEVICE_ID=1003
MM919 331 136 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8232 $Y=1600  $PIN_XY=8262,1594,8232,1600,8202,1594 $DEVICE_ID=1003
MM920 VDD! 136 331 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8064 $Y=1701  $PIN_XY=8094,1594,8064,1701,8034,1594 $DEVICE_ID=1003
MM921 331 136 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7896 $Y=1680  $PIN_XY=7926,1594,7896,1680,7866,1594 $DEVICE_ID=1003
MM922 VDD! 89 135 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7896 $Y=1239  $PIN_XY=7926,1304,7896,1239,7866,1304 $DEVICE_ID=1003
MM923 135 334 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7728 $Y=1218  $PIN_XY=7758,1304,7728,1218,7698,1304 $DEVICE_ID=1003
MM924 VDD! 134 136 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7560 $Y=1600  $PIN_XY=7590,1594,7560,1600,7530,1594 $DEVICE_ID=1003
MM925 136 134 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7392 $Y=1680  $PIN_XY=7422,1594,7392,1680,7362,1594 $DEVICE_ID=1003
MM926 VDD! 92 334 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7392 $Y=1319  $PIN_XY=7422,1304,7392,1319,7362,1304 $DEVICE_ID=1003
MM927 334 92 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7224 $Y=1298  $PIN_XY=7254,1304,7224,1298,7194,1304 $DEVICE_ID=1003
MM928 VDD! D<0> 134 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7056 $Y=1579  $PIN_XY=7086,1594,7056,1579,7026,1594 $DEVICE_ID=1003
MM929 VDD! 92 334 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7056 $Y=1239  $PIN_XY=7086,1304,7056,1239,7026,1304 $DEVICE_ID=1003
MM930 134 D<0> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=1680  $PIN_XY=6918,1594,6888,1680,6858,1594 $DEVICE_ID=1003
MM931 334 92 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6888 $Y=1239  $PIN_XY=6918,1304,6888,1239,6858,1304 $DEVICE_ID=1003
MM932 VDD! 106 107 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6552 $Y=1298  $PIN_XY=6582,1304,6552,1298,6522,1304 $DEVICE_ID=1003
MM933 107 106 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6384 $Y=1218  $PIN_XY=6414,1304,6384,1218,6354,1304 $DEVICE_ID=1003
MM934 VDD! WENB 106 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5880 $Y=1218  $PIN_XY=5910,1304,5880,1218,5850,1304 $DEVICE_ID=1003
MM935 106 102 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5712 $Y=1218  $PIN_XY=5742,1304,5712,1218,5682,1304 $DEVICE_ID=1003
MM936 VDD! 307 78 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5376 $Y=676  $PIN_XY=5406,670,5376,676,5346,670 $DEVICE_ID=1003
MM937 78 307 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5208 $Y=676  $PIN_XY=5238,670,5208,676,5178,670 $DEVICE_ID=1003
MM938 VDD! 307 78 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5040 $Y=777  $PIN_XY=5070,670,5040,777,5010,670 $DEVICE_ID=1003
MM939 78 307 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4872 $Y=777  $PIN_XY=4902,670,4872,777,4842,670 $DEVICE_ID=1003
MM940 VDD! 510 306 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4536 $Y=777  $PIN_XY=4566,670,4536,777,4506,670 $DEVICE_ID=1003
MM941 306 509 307 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4368 $Y=777  $PIN_XY=4398,670,4368,777,4338,670 $DEVICE_ID=1003
XXB19A871F1 GND! VDD! 107 106 274 294 inv $T=6162 924 0 0 $X=6162 $Y=924
XXB19A871F2 VDD! GND! VDD! D<0> 136 332 91 88 134 333 92 
+	92 92 135 _GENERATED_550 _GENERATED_552 _GENERATED_551 _GENERATED_553 89 276 294 295 
+	331 Write_Driver $T=6518 828 0 0 $X=6665 $Y=1384
XXB19A871F3 VDD! GND! VDD! D<1> 139 336 95 93 137 337 96 
+	96 96 138 _GENERATED_554 _GENERATED_556 _GENERATED_555 _GENERATED_557 94 276 294 295 
+	335 Write_Driver $T=9542 828 0 0 $X=9690 $Y=1384
XXB19A871F4 VDD! GND! VDD! D<2> 142 339 86 84 140 340 87 
+	87 87 141 _GENERATED_558 _GENERATED_560 _GENERATED_559 _GENERATED_561 85 276 294 295 
+	338 Write_Driver $T=12566 828 0 0 $X=12714 $Y=1384
XXB19A871F5 VDD! GND! VDD! D<3> 145 342 82 80 143 343 83 
+	83 83 144 VDD! GND! VDD! GND! 81 276 294 295 
+	341 Write_Driver $T=15590 828 0 0 $X=15738 $Y=1384
XXB19A871F6 VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! 310 510 
+	305 WENB 509 308 104 78 77 73 74 103 79 
+	WS0BAR 307 A<1> A<0> 274 275 276 277 294 295 293 
+	292 291 306 309 311 agen_unit $T=1288 2074 0 0 $X=1290 $Y=459
XXB19A871F7 VDD! GND! 8 9 75 146 146 279 15 precharge_logic $T=9462 7518 0 180 $X=8682 $Y=6930
XXB19A871F8 VDD! GND! 10 11 75 147 147 279 15 precharge_logic $T=8790 7518 0 180 $X=8010 $Y=6930
XXB19A871F9 VDD! GND! 12 13 75 148 148 279 15 precharge_logic $T=8118 7518 0 180 $X=7338 $Y=6930
XXB19A871F10 VDD! GND! 14 15 75 149 149 279 15 precharge_logic $T=7446 7518 0 180 $X=6665 $Y=6930
XXB19A871F11 VDD! GND! 23 22 75 158 158 279 15 precharge_logic $T=12486 7518 0 180 $X=11706 $Y=6930
XXB19A871F12 VDD! GND! 21 20 75 159 159 279 15 precharge_logic $T=11814 7518 0 180 $X=11034 $Y=6930
XXB19A871F13 VDD! GND! 19 18 75 160 160 279 15 precharge_logic $T=11142 7518 0 180 $X=10362 $Y=6930
XXB19A871F14 VDD! GND! 16 17 75 161 161 279 15 precharge_logic $T=10470 7518 0 180 $X=9690 $Y=6930
XXB19A871F15 VDD! GND! 32 33 75 182 182 279 15 precharge_logic $T=16518 7518 0 180 $X=15738 $Y=6930
XXB19A871F16 VDD! GND! 34 35 75 183 183 279 15 precharge_logic $T=17190 7518 0 180 $X=16410 $Y=6930
XXB19A871F17 VDD! GND! 36 37 75 184 184 279 15 precharge_logic $T=17862 7518 0 180 $X=17082 $Y=6930
XXB19A871F18 VDD! GND! 38 39 75 185 185 279 15 precharge_logic $T=18534 7518 0 180 $X=17753 $Y=6930
XXB19A871F19 VDD! GND! 31 30 75 170 170 279 15 precharge_logic $T=15510 7518 0 180 $X=14730 $Y=6930
XXB19A871F20 VDD! GND! 24 25 75 171 171 279 15 precharge_logic $T=14838 7518 0 180 $X=14058 $Y=6930
XXB19A871F21 VDD! GND! 26 27 75 172 172 279 15 precharge_logic $T=14166 7518 0 180 $X=13386 $Y=6930
XXB19A871F22 VDD! GND! 28 29 75 173 173 279 15 precharge_logic $T=13494 7518 0 180 $X=12714 $Y=6930
XXB19A871F23 GND! VDD! 106 102 WENB 485 274 294 nand $T=5072 696 0 0 $X=5490 $Y=924
XXB19A871F24 GND! VDD! VDD! GND! VDD! GND! VDD! GND! VDD! 313 314 
+	114 113 77 78 103 79 WS0BAR 73 104 76 100 
+	101 98 74 97 108 90 117 277 278 280 281 
+	292 291 296 15 15 312 between_blocks $T=5162 4502 0 0 $X=5490 $Y=3231
XXB19A871F25 GND! VDD! GND! VDD! VDD! GND! GND! 511 479 512 481 
+	513 516 CLK 483 477 102 475 515 113 114 75 
+	478 480 482 484 279 281 280 278 15 296 15 
+	476 WLRef_PC $T=-394 4618 0 0 $X=-53 $Y=4620
XXB19A871F26 GND! VDD! _GENERATED_563 _GENERATED_562 59 60 288 302 Filler $T=-58 14910 1 0 $X=-54 $Y=14320
XXB19A871F27 GND! VDD! _GENERATED_565 _GENERATED_564 61 62 287 302 Filler $T=-58 13860 0 0 $X=-54 $Y=13860
XXB19A871F28 GND! VDD! _GENERATED_567 _GENERATED_566 63 64 287 303 Filler $T=-58 13986 1 0 $X=-54 $Y=13396
XXB19A871F29 GND! VDD! _GENERATED_569 _GENERATED_568 65 66 286 303 Filler $T=-58 12936 0 0 $X=-54 $Y=12936
XXB19A871F30 GND! VDD! _GENERATED_571 _GENERATED_570 67 68 285 304 Filler $T=-58 12012 0 0 $X=-54 $Y=12012
XXB19A871F31 GND! VDD! _GENERATED_573 _GENERATED_572 69 70 286 304 Filler $T=-58 13062 1 0 $X=-54 $Y=12472
XXB19A871F32 GND! VDD! _GENERATED_575 _GENERATED_574 43 44 284 300 Filler $T=-58 11088 0 0 $X=-54 $Y=11088
XXB19A871F33 GND! VDD! _GENERATED_577 _GENERATED_576 71 72 285 300 Filler $T=-58 12138 1 0 $X=-54 $Y=11548
XXB19A871F34 GND! VDD! _GENERATED_579 _GENERATED_578 45 46 284 301 Filler $T=-58 11214 1 0 $X=-54 $Y=10624
XXB19A871F35 GND! VDD! _GENERATED_581 _GENERATED_580 47 48 283 301 Filler $T=-58 10164 0 0 $X=-54 $Y=10164
XXB19A871F36 GND! VDD! _GENERATED_583 _GENERATED_582 49 50 283 299 Filler $T=-58 10290 1 0 $X=-54 $Y=9700
XXB19A871F37 GND! VDD! _GENERATED_585 _GENERATED_584 51 52 282 299 Filler $T=-58 9240 0 0 $X=-54 $Y=9240
XXB19A871F38 GND! VDD! _GENERATED_587 _GENERATED_586 53 54 282 297 Filler $T=-58 9366 1 0 $X=-54 $Y=8776
XXB19A871F39 GND! VDD! _GENERATED_589 _GENERATED_588 55 56 289 297 Filler $T=-58 8316 0 0 $X=-54 $Y=8316
XXB19A871F40 GND! VDD! _GENERATED_591 _GENERATED_590 57 58 289 298 Filler $T=-58 8442 1 0 $X=-54 $Y=7852
XXB19A871F41 GND! VDD! _GENERATED_593 _GENERATED_592 41 42 279 298 Filler $T=-58 7392 0 0 $X=-54 $Y=7392
XXB19A871F42 GND! VDD! 59 60 _GENERATED_595 _GENERATED_594 288 302 Filler $T=110 14910 1 0 $X=114 $Y=14320
XXB19A871F43 GND! VDD! 61 62 _GENERATED_597 _GENERATED_596 287 302 Filler $T=110 13860 0 0 $X=114 $Y=13860
XXB19A871F44 GND! VDD! 63 64 _GENERATED_599 _GENERATED_598 287 303 Filler $T=110 13986 1 0 $X=114 $Y=13396
XXB19A871F45 GND! VDD! 65 66 _GENERATED_601 _GENERATED_600 286 303 Filler $T=110 12936 0 0 $X=114 $Y=12936
XXB19A871F46 GND! VDD! 67 68 _GENERATED_603 _GENERATED_602 285 304 Filler $T=110 12012 0 0 $X=114 $Y=12012
XXB19A871F47 GND! VDD! 69 70 _GENERATED_605 _GENERATED_604 286 304 Filler $T=110 13062 1 0 $X=114 $Y=12472
XXB19A871F48 GND! VDD! 43 44 _GENERATED_607 _GENERATED_606 284 300 Filler $T=110 11088 0 0 $X=114 $Y=11088
XXB19A871F49 GND! VDD! 71 72 _GENERATED_609 _GENERATED_608 285 300 Filler $T=110 12138 1 0 $X=114 $Y=11548
XXB19A871F50 GND! VDD! 55 56 _GENERATED_611 _GENERATED_610 289 297 Filler $T=110 8316 0 0 $X=114 $Y=8316
XXB19A871F51 GND! VDD! 41 42 _GENERATED_613 _GENERATED_612 279 298 Filler $T=110 7392 0 0 $X=114 $Y=7392
XXB19A871F52 GND! VDD! 57 58 _GENERATED_615 _GENERATED_614 289 298 Filler $T=110 8442 1 0 $X=114 $Y=7852
XXB19A871F53 GND! VDD! 53 54 _GENERATED_617 _GENERATED_616 282 297 Filler $T=110 9366 1 0 $X=114 $Y=8776
XXB19A871F54 GND! VDD! 45 46 _GENERATED_619 _GENERATED_618 284 301 Filler $T=110 11214 1 0 $X=114 $Y=10624
XXB19A871F55 GND! VDD! 47 48 _GENERATED_621 _GENERATED_620 283 301 Filler $T=110 10164 0 0 $X=114 $Y=10164
XXB19A871F56 GND! VDD! 49 50 _GENERATED_623 _GENERATED_622 283 299 Filler $T=110 10290 1 0 $X=114 $Y=9700
XXB19A871F57 GND! VDD! 51 52 _GENERATED_625 _GENERATED_624 282 299 Filler $T=110 9240 0 0 $X=114 $Y=9240
XXB19A871F58 GND! VDD! _GENERATED_628 _GENERATED_626 _GENERATED_629 _GENERATED_627 279 298 Filler $T=446 7392 0 0 $X=450 $Y=7392
XXB19A871F59 GND! VDD! _GENERATED_632 _GENERATED_630 _GENERATED_633 _GENERATED_631 289 298 Filler $T=446 8442 1 0 $X=450 $Y=7852
XXB19A871F60 GND! VDD! _GENERATED_636 _GENERATED_634 _GENERATED_637 _GENERATED_635 289 297 Filler $T=446 8316 0 0 $X=450 $Y=8316
XXB19A871F61 GND! VDD! _GENERATED_640 _GENERATED_638 _GENERATED_641 _GENERATED_639 282 297 Filler $T=446 9366 1 0 $X=450 $Y=8776
XXB19A871F62 GND! VDD! _GENERATED_644 _GENERATED_642 _GENERATED_645 _GENERATED_643 282 299 Filler $T=446 9240 0 0 $X=450 $Y=9240
XXB19A871F63 GND! VDD! _GENERATED_648 _GENERATED_646 _GENERATED_649 _GENERATED_647 283 299 Filler $T=446 10290 1 0 $X=450 $Y=9700
XXB19A871F64 GND! VDD! _GENERATED_652 _GENERATED_650 _GENERATED_653 _GENERATED_651 283 301 Filler $T=446 10164 0 0 $X=450 $Y=10164
XXB19A871F65 GND! VDD! _GENERATED_656 _GENERATED_654 _GENERATED_657 _GENERATED_655 284 301 Filler $T=446 11214 1 0 $X=450 $Y=10624
XXB19A871F66 GND! VDD! _GENERATED_660 _GENERATED_658 _GENERATED_661 _GENERATED_659 285 300 Filler $T=446 12138 1 0 $X=450 $Y=11548
XXB19A871F67 GND! VDD! _GENERATED_664 _GENERATED_662 _GENERATED_665 _GENERATED_663 284 300 Filler $T=446 11088 0 0 $X=450 $Y=11088
XXB19A871F68 GND! VDD! _GENERATED_668 _GENERATED_666 _GENERATED_669 _GENERATED_667 286 304 Filler $T=446 13062 1 0 $X=450 $Y=12472
XXB19A871F69 GND! VDD! _GENERATED_672 _GENERATED_670 _GENERATED_673 _GENERATED_671 285 304 Filler $T=446 12012 0 0 $X=450 $Y=12012
XXB19A871F70 GND! VDD! _GENERATED_676 _GENERATED_674 _GENERATED_677 _GENERATED_675 286 303 Filler $T=446 12936 0 0 $X=450 $Y=12936
XXB19A871F71 GND! VDD! _GENERATED_680 _GENERATED_678 _GENERATED_681 _GENERATED_679 287 303 Filler $T=446 13986 1 0 $X=450 $Y=13396
XXB19A871F72 GND! VDD! _GENERATED_684 _GENERATED_682 _GENERATED_685 _GENERATED_683 287 302 Filler $T=446 13860 0 0 $X=450 $Y=13860
XXB19A871F73 GND! VDD! _GENERATED_688 _GENERATED_686 _GENERATED_689 _GENERATED_687 288 302 Filler $T=446 14910 1 0 $X=450 $Y=14320
XXB19A871F74 GND! VDD! _GENERATED_692 _GENERATED_690 _GENERATED_693 _GENERATED_691 282 299 Filler $T=782 9240 0 0 $X=786 $Y=9240
XXB19A871F75 GND! VDD! _GENERATED_696 _GENERATED_694 _GENERATED_697 _GENERATED_695 283 299 Filler $T=782 10290 1 0 $X=786 $Y=9700
XXB19A871F76 GND! VDD! _GENERATED_700 _GENERATED_698 _GENERATED_701 _GENERATED_699 283 301 Filler $T=782 10164 0 0 $X=786 $Y=10164
XXB19A871F77 GND! VDD! _GENERATED_704 _GENERATED_702 _GENERATED_705 _GENERATED_703 284 301 Filler $T=782 11214 1 0 $X=786 $Y=10624
XXB19A871F78 GND! VDD! _GENERATED_708 _GENERATED_706 _GENERATED_709 _GENERATED_707 282 297 Filler $T=782 9366 1 0 $X=786 $Y=8776
XXB19A871F79 GND! VDD! _GENERATED_712 _GENERATED_710 _GENERATED_713 _GENERATED_711 289 298 Filler $T=782 8442 1 0 $X=786 $Y=7852
XXB19A871F80 GND! VDD! _GENERATED_716 _GENERATED_714 _GENERATED_717 _GENERATED_715 279 298 Filler $T=782 7392 0 0 $X=786 $Y=7392
XXB19A871F81 GND! VDD! _GENERATED_720 _GENERATED_718 _GENERATED_721 _GENERATED_719 289 297 Filler $T=782 8316 0 0 $X=786 $Y=8316
XXB19A871F82 GND! VDD! _GENERATED_724 _GENERATED_722 _GENERATED_725 _GENERATED_723 285 300 Filler $T=782 12138 1 0 $X=786 $Y=11548
XXB19A871F83 GND! VDD! _GENERATED_728 _GENERATED_726 _GENERATED_729 _GENERATED_727 284 300 Filler $T=782 11088 0 0 $X=786 $Y=11088
XXB19A871F84 GND! VDD! _GENERATED_732 _GENERATED_730 _GENERATED_733 _GENERATED_731 286 304 Filler $T=782 13062 1 0 $X=786 $Y=12472
XXB19A871F85 GND! VDD! _GENERATED_736 _GENERATED_734 _GENERATED_737 _GENERATED_735 285 304 Filler $T=782 12012 0 0 $X=786 $Y=12012
XXB19A871F86 GND! VDD! _GENERATED_740 _GENERATED_738 _GENERATED_741 _GENERATED_739 286 303 Filler $T=782 12936 0 0 $X=786 $Y=12936
XXB19A871F87 GND! VDD! _GENERATED_744 _GENERATED_742 _GENERATED_745 _GENERATED_743 287 303 Filler $T=782 13986 1 0 $X=786 $Y=13396
XXB19A871F88 GND! VDD! _GENERATED_748 _GENERATED_746 _GENERATED_749 _GENERATED_747 287 302 Filler $T=782 13860 0 0 $X=786 $Y=13860
XXB19A871F89 GND! VDD! _GENERATED_752 _GENERATED_750 _GENERATED_753 _GENERATED_751 288 302 Filler $T=782 14910 1 0 $X=786 $Y=14320
XXB19A871F90 GND! VDD! _GENERATED_756 _GENERATED_754 _GENERATED_757 _GENERATED_755 288 302 Filler $T=1118 14910 1 0 $X=1122 $Y=14320
XXB19A871F91 GND! VDD! _GENERATED_760 _GENERATED_758 _GENERATED_761 _GENERATED_759 287 302 Filler $T=1118 13860 0 0 $X=1122 $Y=13860
XXB19A871F92 GND! VDD! _GENERATED_764 _GENERATED_762 _GENERATED_765 _GENERATED_763 287 303 Filler $T=1118 13986 1 0 $X=1122 $Y=13396
XXB19A871F93 GND! VDD! _GENERATED_768 _GENERATED_766 _GENERATED_769 _GENERATED_767 286 303 Filler $T=1118 12936 0 0 $X=1122 $Y=12936
XXB19A871F94 GND! VDD! _GENERATED_772 _GENERATED_770 _GENERATED_773 _GENERATED_771 285 304 Filler $T=1118 12012 0 0 $X=1122 $Y=12012
XXB19A871F95 GND! VDD! _GENERATED_776 _GENERATED_774 _GENERATED_777 _GENERATED_775 286 304 Filler $T=1118 13062 1 0 $X=1122 $Y=12472
XXB19A871F96 GND! VDD! _GENERATED_780 _GENERATED_778 _GENERATED_781 _GENERATED_779 284 300 Filler $T=1118 11088 0 0 $X=1122 $Y=11088
XXB19A871F97 GND! VDD! _GENERATED_784 _GENERATED_782 _GENERATED_785 _GENERATED_783 285 300 Filler $T=1118 12138 1 0 $X=1122 $Y=11548
XXB19A871F98 GND! VDD! _GENERATED_788 _GENERATED_786 _GENERATED_789 _GENERATED_787 284 301 Filler $T=1118 11214 1 0 $X=1122 $Y=10624
XXB19A871F99 GND! VDD! _GENERATED_792 _GENERATED_790 _GENERATED_793 _GENERATED_791 283 301 Filler $T=1118 10164 0 0 $X=1122 $Y=10164
XXB19A871F100 GND! VDD! _GENERATED_796 _GENERATED_794 _GENERATED_797 _GENERATED_795 283 299 Filler $T=1118 10290 1 0 $X=1122 $Y=9700
XXB19A871F101 GND! VDD! _GENERATED_800 _GENERATED_798 _GENERATED_801 _GENERATED_799 282 299 Filler $T=1118 9240 0 0 $X=1122 $Y=9240
XXB19A871F102 GND! VDD! _GENERATED_804 _GENERATED_802 _GENERATED_805 _GENERATED_803 282 297 Filler $T=1118 9366 1 0 $X=1122 $Y=8776
XXB19A871F103 GND! VDD! _GENERATED_808 _GENERATED_806 _GENERATED_809 _GENERATED_807 289 297 Filler $T=1118 8316 0 0 $X=1122 $Y=8316
XXB19A871F104 GND! VDD! _GENERATED_812 _GENERATED_810 _GENERATED_813 _GENERATED_811 289 298 Filler $T=1118 8442 1 0 $X=1122 $Y=7852
XXB19A871F105 GND! VDD! _GENERATED_816 _GENERATED_814 _GENERATED_817 _GENERATED_815 279 298 Filler $T=1118 7392 0 0 $X=1122 $Y=7392
XXB19A871F106 GND! VDD! _GENERATED_820 _GENERATED_818 _GENERATED_821 _GENERATED_819 288 302 Filler $T=1454 14910 1 0 $X=1458 $Y=14320
XXB19A871F107 GND! VDD! _GENERATED_824 _GENERATED_822 _GENERATED_825 _GENERATED_823 287 302 Filler $T=1454 13860 0 0 $X=1458 $Y=13860
XXB19A871F108 GND! VDD! _GENERATED_828 _GENERATED_826 _GENERATED_829 _GENERATED_827 287 303 Filler $T=1454 13986 1 0 $X=1458 $Y=13396
XXB19A871F109 GND! VDD! _GENERATED_832 _GENERATED_830 _GENERATED_833 _GENERATED_831 286 303 Filler $T=1454 12936 0 0 $X=1458 $Y=12936
XXB19A871F110 GND! VDD! _GENERATED_836 _GENERATED_834 _GENERATED_837 _GENERATED_835 285 304 Filler $T=1454 12012 0 0 $X=1458 $Y=12012
XXB19A871F111 GND! VDD! _GENERATED_840 _GENERATED_838 _GENERATED_841 _GENERATED_839 286 304 Filler $T=1454 13062 1 0 $X=1458 $Y=12472
XXB19A871F112 GND! VDD! _GENERATED_844 _GENERATED_842 _GENERATED_845 _GENERATED_843 284 300 Filler $T=1454 11088 0 0 $X=1458 $Y=11088
XXB19A871F113 GND! VDD! _GENERATED_848 _GENERATED_846 _GENERATED_849 _GENERATED_847 285 300 Filler $T=1454 12138 1 0 $X=1458 $Y=11548
XXB19A871F114 GND! VDD! _GENERATED_852 _GENERATED_850 _GENERATED_853 _GENERATED_851 289 297 Filler $T=1454 8316 0 0 $X=1458 $Y=8316
XXB19A871F115 GND! VDD! _GENERATED_856 _GENERATED_854 _GENERATED_857 _GENERATED_855 279 298 Filler $T=1454 7392 0 0 $X=1458 $Y=7392
XXB19A871F116 GND! VDD! _GENERATED_860 _GENERATED_858 _GENERATED_861 _GENERATED_859 289 298 Filler $T=1454 8442 1 0 $X=1458 $Y=7852
XXB19A871F117 GND! VDD! _GENERATED_864 _GENERATED_862 _GENERATED_865 _GENERATED_863 282 297 Filler $T=1454 9366 1 0 $X=1458 $Y=8776
XXB19A871F118 GND! VDD! _GENERATED_868 _GENERATED_866 _GENERATED_869 _GENERATED_867 284 301 Filler $T=1454 11214 1 0 $X=1458 $Y=10624
XXB19A871F119 GND! VDD! _GENERATED_872 _GENERATED_870 _GENERATED_873 _GENERATED_871 283 301 Filler $T=1454 10164 0 0 $X=1458 $Y=10164
XXB19A871F120 GND! VDD! _GENERATED_876 _GENERATED_874 _GENERATED_877 _GENERATED_875 283 299 Filler $T=1454 10290 1 0 $X=1458 $Y=9700
XXB19A871F121 GND! VDD! _GENERATED_880 _GENERATED_878 _GENERATED_881 _GENERATED_879 282 299 Filler $T=1454 9240 0 0 $X=1458 $Y=9240
XXB19A871F122 GND! VDD! _GENERATED_884 _GENERATED_882 _GENERATED_885 _GENERATED_883 279 298 Filler $T=1790 7392 0 0 $X=1794 $Y=7392
XXB19A871F123 GND! VDD! _GENERATED_888 _GENERATED_886 _GENERATED_889 _GENERATED_887 289 298 Filler $T=1790 8442 1 0 $X=1794 $Y=7852
XXB19A871F124 GND! VDD! _GENERATED_892 _GENERATED_890 _GENERATED_893 _GENERATED_891 289 297 Filler $T=1790 8316 0 0 $X=1794 $Y=8316
XXB19A871F125 GND! VDD! _GENERATED_896 _GENERATED_894 _GENERATED_897 _GENERATED_895 282 297 Filler $T=1790 9366 1 0 $X=1794 $Y=8776
XXB19A871F126 GND! VDD! _GENERATED_900 _GENERATED_898 _GENERATED_901 _GENERATED_899 282 299 Filler $T=1790 9240 0 0 $X=1794 $Y=9240
XXB19A871F127 GND! VDD! _GENERATED_904 _GENERATED_902 _GENERATED_905 _GENERATED_903 283 299 Filler $T=1790 10290 1 0 $X=1794 $Y=9700
XXB19A871F128 GND! VDD! _GENERATED_908 _GENERATED_906 _GENERATED_909 _GENERATED_907 283 301 Filler $T=1790 10164 0 0 $X=1794 $Y=10164
XXB19A871F129 GND! VDD! _GENERATED_912 _GENERATED_910 _GENERATED_913 _GENERATED_911 284 301 Filler $T=1790 11214 1 0 $X=1794 $Y=10624
XXB19A871F130 GND! VDD! _GENERATED_916 _GENERATED_914 _GENERATED_917 _GENERATED_915 285 300 Filler $T=1790 12138 1 0 $X=1794 $Y=11548
XXB19A871F131 GND! VDD! _GENERATED_920 _GENERATED_918 _GENERATED_921 _GENERATED_919 284 300 Filler $T=1790 11088 0 0 $X=1794 $Y=11088
XXB19A871F132 GND! VDD! _GENERATED_924 _GENERATED_922 _GENERATED_925 _GENERATED_923 286 304 Filler $T=1790 13062 1 0 $X=1794 $Y=12472
XXB19A871F133 GND! VDD! _GENERATED_928 _GENERATED_926 _GENERATED_929 _GENERATED_927 285 304 Filler $T=1790 12012 0 0 $X=1794 $Y=12012
XXB19A871F134 GND! VDD! _GENERATED_932 _GENERATED_930 _GENERATED_933 _GENERATED_931 286 303 Filler $T=1790 12936 0 0 $X=1794 $Y=12936
XXB19A871F135 GND! VDD! _GENERATED_936 _GENERATED_934 _GENERATED_937 _GENERATED_935 287 303 Filler $T=1790 13986 1 0 $X=1794 $Y=13396
XXB19A871F136 GND! VDD! _GENERATED_940 _GENERATED_938 _GENERATED_941 _GENERATED_939 287 302 Filler $T=1790 13860 0 0 $X=1794 $Y=13860
XXB19A871F137 GND! VDD! _GENERATED_944 _GENERATED_942 _GENERATED_945 _GENERATED_943 288 302 Filler $T=1790 14910 1 0 $X=1794 $Y=14320
XXB19A871F138 GND! VDD! _GENERATED_948 _GENERATED_946 _GENERATED_949 _GENERATED_947 282 299 Filler $T=2126 9240 0 0 $X=2130 $Y=9240
XXB19A871F139 GND! VDD! _GENERATED_952 _GENERATED_950 _GENERATED_953 _GENERATED_951 283 299 Filler $T=2126 10290 1 0 $X=2130 $Y=9700
XXB19A871F140 GND! VDD! _GENERATED_956 _GENERATED_954 _GENERATED_957 _GENERATED_955 283 301 Filler $T=2126 10164 0 0 $X=2130 $Y=10164
XXB19A871F141 GND! VDD! _GENERATED_960 _GENERATED_958 _GENERATED_961 _GENERATED_959 284 301 Filler $T=2126 11214 1 0 $X=2130 $Y=10624
XXB19A871F142 GND! VDD! _GENERATED_964 _GENERATED_962 _GENERATED_965 _GENERATED_963 282 297 Filler $T=2126 9366 1 0 $X=2130 $Y=8776
XXB19A871F143 GND! VDD! _GENERATED_968 _GENERATED_966 _GENERATED_969 _GENERATED_967 289 298 Filler $T=2126 8442 1 0 $X=2130 $Y=7852
XXB19A871F144 GND! VDD! _GENERATED_972 _GENERATED_970 _GENERATED_973 _GENERATED_971 279 298 Filler $T=2126 7392 0 0 $X=2130 $Y=7392
XXB19A871F145 GND! VDD! _GENERATED_976 _GENERATED_974 _GENERATED_977 _GENERATED_975 289 297 Filler $T=2126 8316 0 0 $X=2130 $Y=8316
XXB19A871F146 GND! VDD! _GENERATED_980 _GENERATED_978 _GENERATED_981 _GENERATED_979 285 300 Filler $T=2126 12138 1 0 $X=2130 $Y=11548
XXB19A871F147 GND! VDD! _GENERATED_984 _GENERATED_982 _GENERATED_985 _GENERATED_983 284 300 Filler $T=2126 11088 0 0 $X=2130 $Y=11088
XXB19A871F148 GND! VDD! _GENERATED_988 _GENERATED_986 _GENERATED_989 _GENERATED_987 286 304 Filler $T=2126 13062 1 0 $X=2130 $Y=12472
XXB19A871F149 GND! VDD! _GENERATED_992 _GENERATED_990 _GENERATED_993 _GENERATED_991 285 304 Filler $T=2126 12012 0 0 $X=2130 $Y=12012
XXB19A871F150 GND! VDD! _GENERATED_996 _GENERATED_994 _GENERATED_997 _GENERATED_995 286 303 Filler $T=2126 12936 0 0 $X=2130 $Y=12936
XXB19A871F151 GND! VDD! _GENERATED_1000 _GENERATED_998 _GENERATED_1001 _GENERATED_999 287 303 Filler $T=2126 13986 1 0 $X=2130 $Y=13396
XXB19A871F152 GND! VDD! _GENERATED_1004 _GENERATED_1002 _GENERATED_1005 _GENERATED_1003 287 302 Filler $T=2126 13860 0 0 $X=2130 $Y=13860
XXB19A871F153 GND! VDD! _GENERATED_1008 _GENERATED_1006 _GENERATED_1009 _GENERATED_1007 288 302 Filler $T=2126 14910 1 0 $X=2130 $Y=14320
XXB19A871F154 GND! VDD! _GENERATED_1012 _GENERATED_1010 _GENERATED_1013 _GENERATED_1011 288 302 Filler $T=2462 14910 1 0 $X=2466 $Y=14320
XXB19A871F155 GND! VDD! _GENERATED_1016 _GENERATED_1014 _GENERATED_1017 _GENERATED_1015 287 302 Filler $T=2462 13860 0 0 $X=2466 $Y=13860
XXB19A871F156 GND! VDD! _GENERATED_1020 _GENERATED_1018 _GENERATED_1021 _GENERATED_1019 287 303 Filler $T=2462 13986 1 0 $X=2466 $Y=13396
XXB19A871F157 GND! VDD! _GENERATED_1024 _GENERATED_1022 _GENERATED_1025 _GENERATED_1023 286 303 Filler $T=2462 12936 0 0 $X=2466 $Y=12936
XXB19A871F158 GND! VDD! _GENERATED_1028 _GENERATED_1026 _GENERATED_1029 _GENERATED_1027 285 304 Filler $T=2462 12012 0 0 $X=2466 $Y=12012
XXB19A871F159 GND! VDD! _GENERATED_1032 _GENERATED_1030 _GENERATED_1033 _GENERATED_1031 286 304 Filler $T=2462 13062 1 0 $X=2466 $Y=12472
XXB19A871F160 GND! VDD! _GENERATED_1036 _GENERATED_1034 _GENERATED_1037 _GENERATED_1035 284 300 Filler $T=2462 11088 0 0 $X=2466 $Y=11088
XXB19A871F161 GND! VDD! _GENERATED_1040 _GENERATED_1038 _GENERATED_1041 _GENERATED_1039 285 300 Filler $T=2462 12138 1 0 $X=2466 $Y=11548
XXB19A871F162 GND! VDD! _GENERATED_1044 _GENERATED_1042 _GENERATED_1045 _GENERATED_1043 284 301 Filler $T=2462 11214 1 0 $X=2466 $Y=10624
XXB19A871F163 GND! VDD! _GENERATED_1048 _GENERATED_1046 _GENERATED_1049 _GENERATED_1047 283 301 Filler $T=2462 10164 0 0 $X=2466 $Y=10164
XXB19A871F164 GND! VDD! _GENERATED_1052 _GENERATED_1050 _GENERATED_1053 _GENERATED_1051 283 299 Filler $T=2462 10290 1 0 $X=2466 $Y=9700
XXB19A871F165 GND! VDD! _GENERATED_1056 _GENERATED_1054 _GENERATED_1057 _GENERATED_1055 282 299 Filler $T=2462 9240 0 0 $X=2466 $Y=9240
XXB19A871F166 GND! VDD! _GENERATED_1060 _GENERATED_1058 _GENERATED_1061 _GENERATED_1059 282 297 Filler $T=2462 9366 1 0 $X=2466 $Y=8776
XXB19A871F167 GND! VDD! _GENERATED_1064 _GENERATED_1062 _GENERATED_1065 _GENERATED_1063 289 297 Filler $T=2462 8316 0 0 $X=2466 $Y=8316
XXB19A871F168 GND! VDD! _GENERATED_1068 _GENERATED_1066 _GENERATED_1069 _GENERATED_1067 289 298 Filler $T=2462 8442 1 0 $X=2466 $Y=7852
XXB19A871F169 GND! VDD! _GENERATED_1072 _GENERATED_1070 _GENERATED_1073 _GENERATED_1071 279 298 Filler $T=2462 7392 0 0 $X=2466 $Y=7392
XXB19A871F170 GND! VDD! _GENERATED_1076 _GENERATED_1074 _GENERATED_1077 _GENERATED_1075 288 302 Filler $T=2798 14910 1 0 $X=2802 $Y=14320
XXB19A871F171 GND! VDD! _GENERATED_1080 _GENERATED_1078 _GENERATED_1081 _GENERATED_1079 287 302 Filler $T=2798 13860 0 0 $X=2802 $Y=13860
XXB19A871F172 GND! VDD! _GENERATED_1084 _GENERATED_1082 _GENERATED_1085 _GENERATED_1083 287 303 Filler $T=2798 13986 1 0 $X=2802 $Y=13396
XXB19A871F173 GND! VDD! _GENERATED_1088 _GENERATED_1086 _GENERATED_1089 _GENERATED_1087 286 303 Filler $T=2798 12936 0 0 $X=2802 $Y=12936
XXB19A871F174 GND! VDD! _GENERATED_1092 _GENERATED_1090 _GENERATED_1093 _GENERATED_1091 285 304 Filler $T=2798 12012 0 0 $X=2802 $Y=12012
XXB19A871F175 GND! VDD! _GENERATED_1096 _GENERATED_1094 _GENERATED_1097 _GENERATED_1095 286 304 Filler $T=2798 13062 1 0 $X=2802 $Y=12472
XXB19A871F176 GND! VDD! _GENERATED_1100 _GENERATED_1098 _GENERATED_1101 _GENERATED_1099 284 300 Filler $T=2798 11088 0 0 $X=2802 $Y=11088
XXB19A871F177 GND! VDD! _GENERATED_1104 _GENERATED_1102 _GENERATED_1105 _GENERATED_1103 285 300 Filler $T=2798 12138 1 0 $X=2802 $Y=11548
XXB19A871F178 GND! VDD! _GENERATED_1108 _GENERATED_1106 _GENERATED_1109 _GENERATED_1107 289 297 Filler $T=2798 8316 0 0 $X=2802 $Y=8316
XXB19A871F179 GND! VDD! _GENERATED_1112 _GENERATED_1110 _GENERATED_1113 _GENERATED_1111 279 298 Filler $T=2798 7392 0 0 $X=2802 $Y=7392
XXB19A871F180 GND! VDD! _GENERATED_1116 _GENERATED_1114 _GENERATED_1117 _GENERATED_1115 289 298 Filler $T=2798 8442 1 0 $X=2802 $Y=7852
XXB19A871F181 GND! VDD! _GENERATED_1120 _GENERATED_1118 _GENERATED_1121 _GENERATED_1119 282 297 Filler $T=2798 9366 1 0 $X=2802 $Y=8776
XXB19A871F182 GND! VDD! _GENERATED_1124 _GENERATED_1122 _GENERATED_1125 _GENERATED_1123 284 301 Filler $T=2798 11214 1 0 $X=2802 $Y=10624
XXB19A871F183 GND! VDD! _GENERATED_1128 _GENERATED_1126 _GENERATED_1129 _GENERATED_1127 283 301 Filler $T=2798 10164 0 0 $X=2802 $Y=10164
XXB19A871F184 GND! VDD! _GENERATED_1132 _GENERATED_1130 _GENERATED_1133 _GENERATED_1131 283 299 Filler $T=2798 10290 1 0 $X=2802 $Y=9700
XXB19A871F185 GND! VDD! _GENERATED_1136 _GENERATED_1134 _GENERATED_1137 _GENERATED_1135 282 299 Filler $T=2798 9240 0 0 $X=2802 $Y=9240
XXB19A871F186 GND! VDD! _GENERATED_1138 VDD! GND! 40 275 295 Filler $T=18874 2898 0 180 $X=18426 $Y=2308
XXB19A871F187 GND! VDD! GND! _GENERATED_1139 _GENERATED_1140 VDD! 275 292 Filler $T=18422 2772 0 0 $X=18426 $Y=2772
XXB19A871F188 GND! VDD! GND! _GENERATED_1141 _GENERATED_1142 VDD! 281 15 Filler $T=18422 6468 0 0 $X=18426 $Y=6468
XXB19A871F189 GND! VDD! _GENERATED_1144 VDD! GND! _GENERATED_1143 281 15 Filler $T=18874 6594 0 180 $X=18426 $Y=6004
XXB19A871F190 GND! VDD! GND! _GENERATED_1145 _GENERATED_1146 VDD! 280 15 Filler $T=18422 5544 0 0 $X=18426 $Y=5544
XXB19A871F191 GND! VDD! _GENERATED_1148 VDD! GND! _GENERATED_1147 280 296 Filler $T=18874 5670 0 180 $X=18426 $Y=5080
XXB19A871F192 GND! VDD! GND! _GENERATED_1149 _GENERATED_1150 VDD! 277 291 Filler $T=18422 3696 0 0 $X=18426 $Y=3696
XXB19A871F193 GND! VDD! _GENERATED_1152 VDD! GND! _GENERATED_1151 277 292 Filler $T=18874 3822 0 180 $X=18426 $Y=3232
XXB19A871F194 GND! VDD! _GENERATED_1154 VDD! GND! _GENERATED_1153 278 291 Filler $T=18874 4746 0 180 $X=18426 $Y=4156
XXB19A871F195 GND! VDD! GND! _GENERATED_1155 _GENERATED_1156 VDD! 278 296 Filler $T=18422 4620 0 0 $X=18426 $Y=4620
XXB19A871F196 GND! VDD! _GENERATED_1159 _GENERATED_1157 _GENERATED_1160 _GENERATED_1158 279 15 Filler $T=9802 7518 0 180 $X=9354 $Y=6928
XXB19A871F197 GND! VDD! _GENERATED_1163 _GENERATED_1161 _GENERATED_1164 _GENERATED_1162 279 15 Filler $T=12826 7518 0 180 $X=12378 $Y=6928
XXB19A871F198 GND! VDD! _GENERATED_1167 _GENERATED_1165 _GENERATED_1168 _GENERATED_1166 279 15 Filler $T=15850 7518 0 180 $X=15402 $Y=6928
XXB19A871F199 GND! VDD! _GENERATED_1170 VDD! GND! _GENERATED_1169 279 15 Filler $T=18874 7518 0 180 $X=18426 $Y=6928
XXB19A871F200 GND! VDD! Q<3> 112 107 290 274 293 tspc_pos_ff $T=17136 0 1 180 $X=15738 $Y=0
XXB19A871F201 GND! VDD! Q<2> 111 107 290 274 293 tspc_pos_ff $T=14112 0 1 180 $X=12714 $Y=0
XXB19A871F202 GND! VDD! Q<1> 110 107 290 274 293 tspc_pos_ff $T=11088 0 1 180 $X=9690 $Y=0
XXB19A871F203 GND! VDD! Q<0> 109 107 290 274 293 tspc_pos_ff $T=8064 0 1 180 $X=6666 $Y=0
XXB19A871F204 VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! 33 32 
+	35 34 37 36 39 38 80 81 82 83 100 
+	90 108 98 182 183 184 185 101 76 315 117 
+	97 316 317 318 278 277 280 281 296 291 292 
+	15 15 2to4_decoder_static $T=15738 3234 0 0 $X=15738 $Y=3232
XXB19A871F205 VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! 29 28 
+	27 26 25 24 30 31 84 85 86 87 100 
+	90 108 98 173 172 171 170 101 76 319 117 
+	97 320 321 322 278 277 280 281 296 291 292 
+	15 15 2to4_decoder_static $T=12714 3234 0 0 $X=12714 $Y=3232
XXB19A871F206 VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! 15 14 
+	13 12 11 10 9 8 88 89 91 92 100 
+	90 108 98 149 148 147 146 101 76 323 117 
+	97 324 325 326 278 277 280 281 296 291 292 
+	15 15 2to4_decoder_static $T=6666 3234 0 0 $X=6666 $Y=3232
XXB19A871F207 VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! 17 16 
+	18 19 20 21 22 23 93 94 95 96 100 
+	90 108 98 161 160 159 158 101 76 327 117 
+	97 328 329 330 278 277 280 281 296 291 292 
+	15 15 2to4_decoder_static $T=9690 3234 0 0 $X=9690 $Y=3232
XXB19A871F208 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=8508 7392 0 0 $X=8508 $Y=7392
XXB19A871F209 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=7836 7392 0 0 $X=7836 $Y=7392
XXB19A871F210 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=7164 7392 0 0 $X=7164 $Y=7392
XXB19A871F211 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=7164 8316 0 0 $X=7164 $Y=8316
XXB19A871F212 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=7836 8316 0 0 $X=7836 $Y=8316
XXB19A871F213 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=8508 8316 0 0 $X=8508 $Y=8316
XXB19A871F214 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=9180 8316 0 0 $X=9180 $Y=8316
XXB19A871F215 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=9180 7392 0 0 $X=9180 $Y=7392
XXB19A871F216 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=9180 9240 0 0 $X=9180 $Y=9240
XXB19A871F217 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=7164 9240 0 0 $X=7164 $Y=9240
XXB19A871F218 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=7836 9240 0 0 $X=7836 $Y=9240
XXB19A871F219 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=8508 9240 0 0 $X=8508 $Y=9240
XXB19A871F220 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=9180 10164 0 0 $X=9180 $Y=10164
XXB19A871F221 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=8508 10164 0 0 $X=8508 $Y=10164
XXB19A871F222 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=7836 10164 0 0 $X=7836 $Y=10164
XXB19A871F223 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=7164 10164 0 0 $X=7164 $Y=10164
XXB19A871F224 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=8508 11088 0 0 $X=8508 $Y=11088
XXB19A871F225 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=7836 11088 0 0 $X=7836 $Y=11088
XXB19A871F226 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=7164 11088 0 0 $X=7164 $Y=11088
XXB19A871F227 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=9180 11088 0 0 $X=9180 $Y=11088
XXB19A871F228 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=7164 12012 0 0 $X=7164 $Y=12012
XXB19A871F229 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=7836 12012 0 0 $X=7836 $Y=12012
XXB19A871F230 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=8508 12012 0 0 $X=8508 $Y=12012
XXB19A871F231 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=9180 12012 0 0 $X=9180 $Y=12012
XXB19A871F232 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=9180 12936 0 0 $X=9180 $Y=12936
XXB19A871F233 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=7164 12936 0 0 $X=7164 $Y=12936
XXB19A871F234 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=7836 12936 0 0 $X=7836 $Y=12936
XXB19A871F235 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=8508 12936 0 0 $X=8508 $Y=12936
XXB19A871F236 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=9180 13860 0 0 $X=9180 $Y=13860
XXB19A871F237 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=8508 13860 0 0 $X=8508 $Y=13860
XXB19A871F238 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=7836 13860 0 0 $X=7836 $Y=13860
XXB19A871F239 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=7164 13860 0 0 $X=7164 $Y=13860
XXB19A871F240 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=10188 13860 0 0 $X=10188 $Y=13860
XXB19A871F241 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=10860 13860 0 0 $X=10860 $Y=13860
XXB19A871F242 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=11532 13860 0 0 $X=11532 $Y=13860
XXB19A871F243 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=12204 13860 0 0 $X=12204 $Y=13860
XXB19A871F244 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=11532 12936 0 0 $X=11532 $Y=12936
XXB19A871F245 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=10860 12936 0 0 $X=10860 $Y=12936
XXB19A871F246 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=10188 12936 0 0 $X=10188 $Y=12936
XXB19A871F247 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=12204 12936 0 0 $X=12204 $Y=12936
XXB19A871F248 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=12204 12012 0 0 $X=12204 $Y=12012
XXB19A871F249 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=11532 12012 0 0 $X=11532 $Y=12012
XXB19A871F250 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=10860 12012 0 0 $X=10860 $Y=12012
XXB19A871F251 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=10188 12012 0 0 $X=10188 $Y=12012
XXB19A871F252 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=12204 11088 0 0 $X=12204 $Y=11088
XXB19A871F253 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=10188 11088 0 0 $X=10188 $Y=11088
XXB19A871F254 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=10860 11088 0 0 $X=10860 $Y=11088
XXB19A871F255 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=11532 11088 0 0 $X=11532 $Y=11088
XXB19A871F256 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=10188 10164 0 0 $X=10188 $Y=10164
XXB19A871F257 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=10860 10164 0 0 $X=10860 $Y=10164
XXB19A871F258 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=11532 10164 0 0 $X=11532 $Y=10164
XXB19A871F259 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=12204 10164 0 0 $X=12204 $Y=10164
XXB19A871F260 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=11532 9240 0 0 $X=11532 $Y=9240
XXB19A871F261 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=10860 9240 0 0 $X=10860 $Y=9240
XXB19A871F262 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=10188 9240 0 0 $X=10188 $Y=9240
XXB19A871F263 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=12204 9240 0 0 $X=12204 $Y=9240
XXB19A871F264 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=10188 8316 0 0 $X=10188 $Y=8316
XXB19A871F265 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=10860 8316 0 0 $X=10860 $Y=8316
XXB19A871F266 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=11532 8316 0 0 $X=11532 $Y=8316
XXB19A871F267 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=12204 8316 0 0 $X=12204 $Y=8316
XXB19A871F268 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=12204 7392 0 0 $X=12204 $Y=7392
XXB19A871F269 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=11532 7392 0 0 $X=11532 $Y=7392
XXB19A871F270 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=10188 7392 0 0 $X=10188 $Y=7392
XXB19A871F271 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=10860 7392 0 0 $X=10860 $Y=7392
XXB19A871F272 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=18252 9240 0 0 $X=18252 $Y=9240
XXB19A871F273 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=16236 9240 0 0 $X=16236 $Y=9240
XXB19A871F274 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=16908 9240 0 0 $X=16908 $Y=9240
XXB19A871F275 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=17580 9240 0 0 $X=17580 $Y=9240
XXB19A871F276 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=18252 10164 0 0 $X=18252 $Y=10164
XXB19A871F277 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=17580 10164 0 0 $X=17580 $Y=10164
XXB19A871F278 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=16908 10164 0 0 $X=16908 $Y=10164
XXB19A871F279 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=16236 10164 0 0 $X=16236 $Y=10164
XXB19A871F280 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=17580 11088 0 0 $X=17580 $Y=11088
XXB19A871F281 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=16908 11088 0 0 $X=16908 $Y=11088
XXB19A871F282 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=16236 11088 0 0 $X=16236 $Y=11088
XXB19A871F283 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=18252 11088 0 0 $X=18252 $Y=11088
XXB19A871F284 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=16236 12012 0 0 $X=16236 $Y=12012
XXB19A871F285 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=16908 12012 0 0 $X=16908 $Y=12012
XXB19A871F286 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=17580 12012 0 0 $X=17580 $Y=12012
XXB19A871F287 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=18252 12012 0 0 $X=18252 $Y=12012
XXB19A871F288 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=18252 12936 0 0 $X=18252 $Y=12936
XXB19A871F289 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=16236 12936 0 0 $X=16236 $Y=12936
XXB19A871F290 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=16908 12936 0 0 $X=16908 $Y=12936
XXB19A871F291 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=17580 12936 0 0 $X=17580 $Y=12936
XXB19A871F292 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=18252 13860 0 0 $X=18252 $Y=13860
XXB19A871F293 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=17580 13860 0 0 $X=17580 $Y=13860
XXB19A871F294 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=16908 13860 0 0 $X=16908 $Y=13860
XXB19A871F295 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=16236 13860 0 0 $X=16236 $Y=13860
XXB19A871F296 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=14556 13860 0 0 $X=14556 $Y=13860
XXB19A871F297 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=15228 13860 0 0 $X=15228 $Y=13860
XXB19A871F298 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=14556 12936 0 0 $X=14556 $Y=12936
XXB19A871F299 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=15228 12936 0 0 $X=15228 $Y=12936
XXB19A871F300 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=15228 12012 0 0 $X=15228 $Y=12012
XXB19A871F301 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=14556 12012 0 0 $X=14556 $Y=12012
XXB19A871F302 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=15228 11088 0 0 $X=15228 $Y=11088
XXB19A871F303 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=14556 11088 0 0 $X=14556 $Y=11088
XXB19A871F304 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=14556 10164 0 0 $X=14556 $Y=10164
XXB19A871F305 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=15228 10164 0 0 $X=15228 $Y=10164
XXB19A871F306 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=14556 9240 0 0 $X=14556 $Y=9240
XXB19A871F307 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=15228 9240 0 0 $X=15228 $Y=9240
XXB19A871F308 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=16908 7392 0 0 $X=16908 $Y=7392
XXB19A871F309 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=16236 7392 0 0 $X=16236 $Y=7392
XXB19A871F310 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=17580 7392 0 0 $X=17580 $Y=7392
XXB19A871F311 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=18252 7392 0 0 $X=18252 $Y=7392
XXB19A871F312 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=18252 8316 0 0 $X=18252 $Y=8316
XXB19A871F313 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=17580 8316 0 0 $X=17580 $Y=8316
XXB19A871F314 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=16908 8316 0 0 $X=16908 $Y=8316
XXB19A871F315 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=16236 8316 0 0 $X=16236 $Y=8316
XXB19A871F316 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=13212 13860 0 0 $X=13212 $Y=13860
XXB19A871F317 GND! VDD! GND! 287 288 302 bitcell_precharge_filler $T=13884 13860 0 0 $X=13884 $Y=13860
XXB19A871F318 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=13884 12936 0 0 $X=13884 $Y=12936
XXB19A871F319 GND! VDD! GND! 286 287 303 bitcell_precharge_filler $T=13212 12936 0 0 $X=13212 $Y=12936
XXB19A871F320 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=13884 12012 0 0 $X=13884 $Y=12012
XXB19A871F321 GND! VDD! GND! 285 286 304 bitcell_precharge_filler $T=13212 12012 0 0 $X=13212 $Y=12012
XXB19A871F322 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=13212 11088 0 0 $X=13212 $Y=11088
XXB19A871F323 GND! VDD! GND! 284 285 300 bitcell_precharge_filler $T=13884 11088 0 0 $X=13884 $Y=11088
XXB19A871F324 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=13212 10164 0 0 $X=13212 $Y=10164
XXB19A871F325 GND! VDD! GND! 283 284 301 bitcell_precharge_filler $T=13884 10164 0 0 $X=13884 $Y=10164
XXB19A871F326 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=13884 9240 0 0 $X=13884 $Y=9240
XXB19A871F327 GND! VDD! GND! 282 283 299 bitcell_precharge_filler $T=13212 9240 0 0 $X=13212 $Y=9240
XXB19A871F328 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=13212 8316 0 0 $X=13212 $Y=8316
XXB19A871F329 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=13884 8316 0 0 $X=13884 $Y=8316
XXB19A871F330 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=14556 8316 0 0 $X=14556 $Y=8316
XXB19A871F331 GND! VDD! GND! 289 282 297 bitcell_precharge_filler $T=15228 8316 0 0 $X=15228 $Y=8316
XXB19A871F332 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=15228 7392 0 0 $X=15228 $Y=7392
XXB19A871F333 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=14556 7392 0 0 $X=14556 $Y=7392
XXB19A871F334 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=13212 7392 0 0 $X=13212 $Y=7392
XXB19A871F335 GND! VDD! GND! 279 289 298 bitcell_precharge_filler $T=13884 7392 0 0 $X=13884 $Y=7392
XXB19A871F336 VDD! GND! GND! GND! VDD! VDD! GND! VDD! GND! GND! VDD! 
+	GND! VDD! GND! GND! VDD! 517 A<2> A<3> 514 A<4> 491 
+	113 120 116 121 122 115 119 124 123 279 289 
+	283 282 285 284 288 287 286 298 297 299 301 
+	300 303 304 302 492 490 static_row_decoder_3by8 $T=2486 13270 0 0 $X=3138 $Y=7391
XXB19A871F337 GND! VDD! VDD! GND! 274 293 2to4_decoder_static_filler_17 $T=18870 1054 0 180 $X=18426 $Y=462
XXB19A871F338 GND! VDD! _GENERATED_1172 _GENERATED_1171 274 294 2to4_decoder_static_filler_17 $T=18426 920 0 0 $X=18426 $Y=924
XXB19A871F339 GND! VDD! _GENERATED_1174 _GENERATED_1173 274 294 2to4_decoder_static_filler_17 $T=17754 920 0 0 $X=17754 $Y=924
XXB19A871F340 GND! VDD! _GENERATED_1176 _GENERATED_1175 274 294 2to4_decoder_static_filler_17 $T=18090 920 0 0 $X=18090 $Y=924
XXB19A871F341 GND! VDD! _GENERATED_1178 _GENERATED_1177 274 293 2to4_decoder_static_filler_17 $T=18534 1054 0 180 $X=18090 $Y=462
XXB19A871F342 GND! VDD! _GENERATED_1180 _GENERATED_1179 274 293 2to4_decoder_static_filler_17 $T=18198 1054 0 180 $X=17754 $Y=462
XXB19A871F343 GND! VDD! _GENERATED_1182 _GENERATED_1181 274 293 2to4_decoder_static_filler_17 $T=17526 1054 0 180 $X=17082 $Y=462
XXB19A871F344 GND! VDD! _GENERATED_1184 _GENERATED_1183 274 293 2to4_decoder_static_filler_17 $T=17862 1054 0 180 $X=17418 $Y=462
XXB19A871F345 GND! VDD! _GENERATED_1186 _GENERATED_1185 274 294 2to4_decoder_static_filler_17 $T=14730 920 0 0 $X=14730 $Y=924
XXB19A871F346 GND! VDD! _GENERATED_1188 _GENERATED_1187 274 294 2to4_decoder_static_filler_17 $T=15066 920 0 0 $X=15066 $Y=924
XXB19A871F347 GND! VDD! _GENERATED_1190 _GENERATED_1189 274 294 2to4_decoder_static_filler_17 $T=15402 920 0 0 $X=15402 $Y=924
XXB19A871F348 GND! VDD! _GENERATED_1192 _GENERATED_1191 274 293 2to4_decoder_static_filler_17 $T=15846 1054 0 180 $X=15402 $Y=462
XXB19A871F349 GND! VDD! _GENERATED_1194 _GENERATED_1193 274 293 2to4_decoder_static_filler_17 $T=15510 1054 0 180 $X=15065 $Y=462
XXB19A871F350 GND! VDD! _GENERATED_1196 _GENERATED_1195 274 293 2to4_decoder_static_filler_17 $T=15174 1054 0 180 $X=14729 $Y=462
XXB19A871F351 GND! VDD! _GENERATED_1198 _GENERATED_1197 274 293 2to4_decoder_static_filler_17 $T=14838 1054 0 180 $X=14394 $Y=462
XXB19A871F352 GND! VDD! _GENERATED_1200 _GENERATED_1199 274 293 2to4_decoder_static_filler_17 $T=14502 1054 0 180 $X=14058 $Y=462
XXB19A871F353 GND! VDD! _GENERATED_1202 _GENERATED_1201 274 293 2to4_decoder_static_filler_17 $T=11814 1054 0 180 $X=11370 $Y=462
XXB19A871F354 GND! VDD! _GENERATED_1204 _GENERATED_1203 274 293 2to4_decoder_static_filler_17 $T=11478 1054 0 180 $X=11033 $Y=462
XXB19A871F355 GND! VDD! _GENERATED_1206 _GENERATED_1205 274 293 2to4_decoder_static_filler_17 $T=12150 1054 0 180 $X=11706 $Y=462
XXB19A871F356 GND! VDD! _GENERATED_1208 _GENERATED_1207 274 293 2to4_decoder_static_filler_17 $T=12486 1054 0 180 $X=12042 $Y=462
XXB19A871F357 GND! VDD! _GENERATED_1210 _GENERATED_1209 274 294 2to4_decoder_static_filler_17 $T=12042 920 0 0 $X=12042 $Y=924
XXB19A871F358 GND! VDD! _GENERATED_1212 _GENERATED_1211 274 294 2to4_decoder_static_filler_17 $T=11706 920 0 0 $X=11706 $Y=924
XXB19A871F359 GND! VDD! _GENERATED_1214 _GENERATED_1213 274 294 2to4_decoder_static_filler_17 $T=12378 920 0 0 $X=12378 $Y=924
XXB19A871F360 GND! VDD! _GENERATED_1216 _GENERATED_1215 274 293 2to4_decoder_static_filler_17 $T=12822 1054 0 180 $X=12378 $Y=462
XXB19A871F361 GND! VDD! _GENERATED_1218 _GENERATED_1217 274 293 2to4_decoder_static_filler_17 $T=8454 1054 0 180 $X=8010 $Y=462
XXB19A871F362 GND! VDD! _GENERATED_1220 _GENERATED_1219 274 293 2to4_decoder_static_filler_17 $T=8790 1054 0 180 $X=8346 $Y=462
XXB19A871F363 GND! VDD! _GENERATED_1222 _GENERATED_1221 274 293 2to4_decoder_static_filler_17 $T=9126 1054 0 180 $X=8681 $Y=462
XXB19A871F364 GND! VDD! _GENERATED_1224 _GENERATED_1223 274 293 2to4_decoder_static_filler_17 $T=9462 1054 0 180 $X=9017 $Y=462
XXB19A871F365 GND! VDD! _GENERATED_1226 _GENERATED_1225 274 293 2to4_decoder_static_filler_17 $T=9798 1054 0 180 $X=9354 $Y=462
XXB19A871F366 GND! VDD! _GENERATED_1228 _GENERATED_1227 274 294 2to4_decoder_static_filler_17 $T=9354 920 0 0 $X=9354 $Y=924
XXB19A871F367 GND! VDD! _GENERATED_1230 _GENERATED_1229 274 294 2to4_decoder_static_filler_17 $T=9018 920 0 0 $X=9018 $Y=924
XXB19A871F368 GND! VDD! _GENERATED_1232 _GENERATED_1231 274 294 2to4_decoder_static_filler_17 $T=8682 920 0 0 $X=8682 $Y=924
XXB19A871F369 GND! VDD! 83 344 81 144 112 D<3> D<3> 143 145 
+	145 274 294 489 read_circuit $T=15738 920 0 0 $X=15738 $Y=924
XXB19A871F370 GND! VDD! 87 345 85 141 111 D<2> D<2> 140 142 
+	142 274 294 487 read_circuit $T=12714 920 0 0 $X=12714 $Y=924
XXB19A871F371 GND! VDD! 96 346 94 138 110 D<1> D<1> 137 139 
+	139 274 294 488 read_circuit $T=9690 920 0 0 $X=9690 $Y=924
XXB19A871F372 GND! VDD! 92 334 89 135 109 D<0> D<0> 134 136 
+	136 274 294 486 read_circuit $T=6666 920 0 0 $X=6666 $Y=924
XXB19A871F373 GND! VDD! _GENERATED_1234 _GENERATED_1233 290 293 sram_filler $T=18422 0 0 0 $X=18426 $Y=0
XXB19A871F374 GND! VDD! _GENERATED_1236 _GENERATED_1235 290 293 sram_filler $T=17078 0 0 0 $X=17082 $Y=0
XXB19A871F375 GND! VDD! _GENERATED_1238 _GENERATED_1237 290 293 sram_filler $T=17414 0 0 0 $X=17418 $Y=0
XXB19A871F376 GND! VDD! _GENERATED_1240 _GENERATED_1239 290 293 sram_filler $T=17750 0 0 0 $X=17754 $Y=0
XXB19A871F377 GND! VDD! _GENERATED_1242 _GENERATED_1241 290 293 sram_filler $T=18086 0 0 0 $X=18090 $Y=0
XXB19A871F378 GND! VDD! _GENERATED_1244 _GENERATED_1243 290 293 sram_filler $T=15398 0 0 0 $X=15402 $Y=0
XXB19A871F379 GND! VDD! _GENERATED_1246 _GENERATED_1245 290 293 sram_filler $T=15062 0 0 0 $X=15066 $Y=0
XXB19A871F380 GND! VDD! _GENERATED_1248 _GENERATED_1247 290 293 sram_filler $T=14726 0 0 0 $X=14730 $Y=0
XXB19A871F381 GND! VDD! _GENERATED_1250 _GENERATED_1249 290 293 sram_filler $T=6326 0 0 0 $X=6330 $Y=0
XXB19A871F382 GND! VDD! _GENERATED_1252 _GENERATED_1251 290 293 sram_filler $T=5990 0 0 0 $X=5994 $Y=0
XXB19A871F383 GND! VDD! _GENERATED_1254 _GENERATED_1253 290 293 sram_filler $T=5654 0 0 0 $X=5657 $Y=0
XXB19A871F384 GND! VDD! _GENERATED_1256 _GENERATED_1255 290 293 sram_filler $T=5318 0 0 0 $X=5322 $Y=0
XXB19A871F385 GND! VDD! _GENERATED_1258 _GENERATED_1257 290 293 sram_filler $T=8006 0 0 0 $X=8010 $Y=0
XXB19A871F386 GND! VDD! _GENERATED_1260 _GENERATED_1259 290 293 sram_filler $T=8342 0 0 0 $X=8346 $Y=0
XXB19A871F387 GND! VDD! _GENERATED_1262 _GENERATED_1261 290 293 sram_filler $T=8678 0 0 0 $X=8682 $Y=0
XXB19A871F388 GND! VDD! _GENERATED_1264 _GENERATED_1263 290 293 sram_filler $T=14054 0 0 0 $X=14058 $Y=0
XXB19A871F389 GND! VDD! _GENERATED_1266 _GENERATED_1265 290 293 sram_filler $T=12038 0 0 0 $X=12042 $Y=0
XXB19A871F390 GND! VDD! _GENERATED_1268 _GENERATED_1267 290 293 sram_filler $T=11702 0 0 0 $X=11706 $Y=0
XXB19A871F391 GND! VDD! _GENERATED_1270 _GENERATED_1269 290 293 sram_filler $T=11366 0 0 0 $X=11370 $Y=0
XXB19A871F392 GND! VDD! _GENERATED_1272 _GENERATED_1271 290 293 sram_filler $T=11030 0 0 0 $X=11033 $Y=0
XXB19A871F393 GND! VDD! _GENERATED_1274 _GENERATED_1273 290 293 sram_filler $T=14390 0 0 0 $X=14394 $Y=0
XXB19A871F394 GND! VDD! _GENERATED_1276 _GENERATED_1275 290 293 sram_filler $T=9014 0 0 0 $X=9017 $Y=0
XXB19A871F395 GND! VDD! _GENERATED_1278 _GENERATED_1277 290 293 sram_filler $T=9350 0 0 0 $X=9354 $Y=0
XXB19A871F396 GND! VDD! _GENERATED_1280 _GENERATED_1279 290 293 sram_filler $T=12374 0 0 0 $X=12378 $Y=0
XXB19A871F397 GND! VDD! _GENERATED_1282 _GENERATED_1281 290 293 sram_filler $T=4982 0 0 0 $X=4986 $Y=0
XXB19A871F398 GND! VDD! _GENERATED_1284 _GENERATED_1283 290 293 sram_filler $T=4646 0 0 0 $X=4649 $Y=0
XXB19A871F399 GND! VDD! _GENERATED_1286 _GENERATED_1285 290 293 sram_filler $T=4310 0 0 0 $X=4314 $Y=0
XXB19A871F400 GND! VDD! _GENERATED_1288 _GENERATED_1287 290 293 sram_filler $T=3974 0 0 0 $X=3978 $Y=0
XXB19A871F401 GND! VDD! _GENERATED_1290 _GENERATED_1289 290 293 sram_filler $T=2630 0 0 0 $X=2634 $Y=0
XXB19A871F402 GND! VDD! _GENERATED_1292 _GENERATED_1291 290 293 sram_filler $T=2966 0 0 0 $X=2970 $Y=0
XXB19A871F403 GND! VDD! _GENERATED_1294 _GENERATED_1293 290 293 sram_filler $T=3302 0 0 0 $X=3306 $Y=0
XXB19A871F404 GND! VDD! _GENERATED_1296 _GENERATED_1295 290 293 sram_filler $T=3638 0 0 0 $X=3642 $Y=0
XXB19A871F405 GND! VDD! _GENERATED_1298 _GENERATED_1297 290 293 sram_filler $T=1286 0 0 0 $X=1290 $Y=0
XXB19A871F406 GND! VDD! _GENERATED_1300 _GENERATED_1299 290 293 sram_filler $T=1622 0 0 0 $X=1626 $Y=0
XXB19A871F407 GND! VDD! _GENERATED_1302 _GENERATED_1301 290 293 sram_filler $T=1958 0 0 0 $X=1962 $Y=0
XXB19A871F408 GND! VDD! _GENERATED_1304 _GENERATED_1303 290 293 sram_filler $T=2294 0 0 0 $X=2298 $Y=0
XXB19A871F409 GND! VDD! _GENERATED_1306 _GENERATED_1305 290 293 sram_filler $T=950 0 0 0 $X=954 $Y=0
XXB19A871F410 GND! VDD! _GENERATED_1308 _GENERATED_1307 290 293 sram_filler $T=614 0 0 0 $X=618 $Y=0
XXB19A871F411 GND! VDD! _GENERATED_1310 _GENERATED_1309 290 293 sram_filler $T=278 0 0 0 $X=282 $Y=0
XXB19A871F412 GND! VDD! _GENERATED_1312 _GENERATED_1311 290 293 sram_filler $T=-58 0 0 0 $X=-54 $Y=0
XXB19A871F413 GND! VDD! _GENERATED_1314 _GENERATED_1313 274 294 sram_filler $T=950 924 0 0 $X=954 $Y=924
XXB19A871F414 GND! VDD! _GENERATED_1316 _GENERATED_1315 274 294 sram_filler $T=614 924 0 0 $X=618 $Y=924
XXB19A871F415 GND! VDD! _GENERATED_1318 _GENERATED_1317 274 294 sram_filler $T=278 924 0 0 $X=282 $Y=924
XXB19A871F416 GND! VDD! _GENERATED_1320 _GENERATED_1319 274 294 sram_filler $T=-58 924 0 0 $X=-54 $Y=924
XXB19A871F417 GND! VDD! _GENERATED_1322 _GENERATED_1321 276 295 sram_filler $T=950 1848 0 0 $X=954 $Y=1848
XXB19A871F418 GND! VDD! _GENERATED_1324 _GENERATED_1323 276 295 sram_filler $T=614 1848 0 0 $X=618 $Y=1848
XXB19A871F419 GND! VDD! _GENERATED_1326 _GENERATED_1325 276 295 sram_filler $T=278 1848 0 0 $X=282 $Y=1848
XXB19A871F420 GND! VDD! _GENERATED_1328 _GENERATED_1327 276 295 sram_filler $T=-58 1848 0 0 $X=-54 $Y=1848
XXB19A871F421 GND! VDD! _GENERATED_1330 _GENERATED_1329 275 292 sram_filler $T=-58 2772 0 0 $X=-54 $Y=2772
XXB19A871F422 GND! VDD! _GENERATED_1332 _GENERATED_1331 275 292 sram_filler $T=278 2772 0 0 $X=282 $Y=2772
XXB19A871F423 GND! VDD! _GENERATED_1334 _GENERATED_1333 275 292 sram_filler $T=614 2772 0 0 $X=618 $Y=2772
XXB19A871F424 GND! VDD! _GENERATED_1336 _GENERATED_1335 275 292 sram_filler $T=950 2772 0 0 $X=954 $Y=2772
XXB19A871F425 GND! VDD! _GENERATED_1338 _GENERATED_1337 277 291 sram_filler $T=-58 3696 0 0 $X=-54 $Y=3696
XXB19A871F426 GND! VDD! _GENERATED_1340 _GENERATED_1339 277 291 sram_filler $T=278 3696 0 0 $X=282 $Y=3696
XXB19A871F427 GND! VDD! _GENERATED_1342 _GENERATED_1341 277 291 sram_filler $T=614 3696 0 0 $X=618 $Y=3696
XXB19A871F428 GND! VDD! _GENERATED_1344 _GENERATED_1343 277 291 sram_filler $T=950 3696 0 0 $X=954 $Y=3696
XXB19A871F429 GND! VDD! VDD! _GENERATED_1345 276 295 sram_filler $T=6326 1848 0 0 $X=6330 $Y=1848
XXB19A871F430 GND! VDD! _GENERATED_1347 _GENERATED_1346 276 295 sram_filler $T=5486 1848 0 0 $X=5489 $Y=1848
XXB19A871F431 GND! VDD! _GENERATED_1349 _GENERATED_1348 276 295 sram_filler $T=5822 1848 0 0 $X=5826 $Y=1848
XXB19A871F432 GND! VDD! _GENERATED_1350 GND! 276 295 sram_filler $T=6158 1848 0 0 $X=6162 $Y=1848
XXB19A871F433 GND! VDD! VDD! _GENERATED_1351 275 292 sram_filler $T=18086 2772 0 0 $X=18090 $Y=2772
XXB19A871F434 GND! VDD! _GENERATED_1353 _GENERATED_1352 275 292 sram_filler $T=17582 2772 0 0 $X=17586 $Y=2772
XXB19A871F435 GND! VDD! _GENERATED_1354 GND! 275 292 sram_filler $T=17918 2772 0 0 $X=17922 $Y=2772
XXB19A871F436 GND! VDD! _GENERATED_1356 _GENERATED_1355 275 292 sram_filler $T=17246 2772 0 0 $X=17250 $Y=2772
XXB19A871F437 GND! VDD! _GENERATED_1358 _GENERATED_1357 275 292 sram_filler $T=16910 2772 0 0 $X=16914 $Y=2772
XXB19A871F438 GND! VDD! _GENERATED_1360 _GENERATED_1359 275 292 sram_filler $T=16238 2772 0 0 $X=16242 $Y=2772
XXB19A871F439 GND! VDD! _GENERATED_1362 _GENERATED_1361 275 292 sram_filler $T=16574 2772 0 0 $X=16578 $Y=2772
XXB19A871F440 GND! VDD! _GENERATED_1364 _GENERATED_1363 275 292 sram_filler $T=13550 2772 0 0 $X=13554 $Y=2772
XXB19A871F441 GND! VDD! _GENERATED_1366 _GENERATED_1365 275 292 sram_filler $T=12878 2772 0 0 $X=12882 $Y=2772
XXB19A871F442 GND! VDD! _GENERATED_1368 _GENERATED_1367 275 292 sram_filler $T=13214 2772 0 0 $X=13218 $Y=2772
XXB19A871F443 GND! VDD! _GENERATED_1370 _GENERATED_1369 275 292 sram_filler $T=12542 2772 0 0 $X=12546 $Y=2772
XXB19A871F444 GND! VDD! _GENERATED_1372 _GENERATED_1371 275 292 sram_filler $T=12206 2772 0 0 $X=12209 $Y=2772
XXB19A871F445 GND! VDD! _GENERATED_1374 _GENERATED_1373 275 292 sram_filler $T=11534 2772 0 0 $X=11538 $Y=2772
XXB19A871F446 GND! VDD! _GENERATED_1376 _GENERATED_1375 275 292 sram_filler $T=11870 2772 0 0 $X=11874 $Y=2772
XXB19A871F447 GND! VDD! _GENERATED_1378 _GENERATED_1377 275 292 sram_filler $T=11198 2772 0 0 $X=11202 $Y=2772
XXB19A871F448 GND! VDD! _GENERATED_1380 _GENERATED_1379 275 292 sram_filler $T=10862 2772 0 0 $X=10866 $Y=2772
XXB19A871F449 GND! VDD! _GENERATED_1382 _GENERATED_1381 275 292 sram_filler $T=15566 2772 0 0 $X=15570 $Y=2772
XXB19A871F450 GND! VDD! _GENERATED_1384 _GENERATED_1383 275 292 sram_filler $T=15902 2772 0 0 $X=15906 $Y=2772
XXB19A871F451 GND! VDD! _GENERATED_1386 _GENERATED_1385 275 292 sram_filler $T=15230 2772 0 0 $X=15234 $Y=2772
XXB19A871F452 GND! VDD! _GENERATED_1388 _GENERATED_1387 275 292 sram_filler $T=14894 2772 0 0 $X=14898 $Y=2772
XXB19A871F453 GND! VDD! _GENERATED_1390 _GENERATED_1389 275 292 sram_filler $T=14222 2772 0 0 $X=14226 $Y=2772
XXB19A871F454 GND! VDD! _GENERATED_1392 _GENERATED_1391 275 292 sram_filler $T=14558 2772 0 0 $X=14562 $Y=2772
XXB19A871F455 GND! VDD! _GENERATED_1394 _GENERATED_1393 275 292 sram_filler $T=13886 2772 0 0 $X=13890 $Y=2772
XXB19A871F456 GND! VDD! _GENERATED_1396 _GENERATED_1395 275 292 sram_filler $T=10190 2772 0 0 $X=10193 $Y=2772
XXB19A871F457 GND! VDD! _GENERATED_1398 _GENERATED_1397 275 292 sram_filler $T=10526 2772 0 0 $X=10530 $Y=2772
XXB19A871F458 GND! VDD! _GENERATED_1400 _GENERATED_1399 275 292 sram_filler $T=9854 2772 0 0 $X=9858 $Y=2772
XXB19A871F459 GND! VDD! _GENERATED_1402 _GENERATED_1401 275 292 sram_filler $T=9518 2772 0 0 $X=9522 $Y=2772
XXB19A871F460 GND! VDD! _GENERATED_1404 _GENERATED_1403 275 292 sram_filler $T=8846 2772 0 0 $X=8850 $Y=2772
XXB19A871F461 GND! VDD! _GENERATED_1406 _GENERATED_1405 275 292 sram_filler $T=9182 2772 0 0 $X=9186 $Y=2772
XXB19A871F462 GND! VDD! _GENERATED_1408 _GENERATED_1407 275 292 sram_filler $T=8510 2772 0 0 $X=8514 $Y=2772
XXB19A871F463 GND! VDD! _GENERATED_1410 _GENERATED_1409 275 292 sram_filler $T=8174 2772 0 0 $X=8177 $Y=2772
XXB19A871F464 GND! VDD! _GENERATED_1412 _GENERATED_1411 275 292 sram_filler $T=7502 2772 0 0 $X=7505 $Y=2772
XXB19A871F465 GND! VDD! _GENERATED_1414 _GENERATED_1413 275 292 sram_filler $T=7838 2772 0 0 $X=7842 $Y=2772
XXB19A871F466 GND! VDD! _GENERATED_1416 _GENERATED_1415 275 292 sram_filler $T=7166 2772 0 0 $X=7170 $Y=2772
XXB19A871F467 GND! VDD! _GENERATED_1418 _GENERATED_1417 275 292 sram_filler $T=6830 2772 0 0 $X=6834 $Y=2772
XXB19A871F468 GND! VDD! _GENERATED_1420 _GENERATED_1419 275 292 sram_filler $T=6158 2772 0 0 $X=6162 $Y=2772
XXB19A871F469 GND! VDD! _GENERATED_1422 _GENERATED_1421 275 292 sram_filler $T=6494 2772 0 0 $X=6497 $Y=2772
XXB19A871F470 GND! VDD! _GENERATED_1424 _GENERATED_1423 275 292 sram_filler $T=5822 2772 0 0 $X=5826 $Y=2772
XXB19A871F471 GND! VDD! _GENERATED_1426 _GENERATED_1425 275 292 sram_filler $T=5486 2772 0 0 $X=5489 $Y=2772
XXB19A871F472 GND! VDD! _GENERATED_1428 _GENERATED_1427 281 15 sram_filler $T=15398 6468 0 0 $X=15402 $Y=6468
XXB19A871F473 GND! VDD! _GENERATED_1430 _GENERATED_1429 280 15 sram_filler $T=15398 5544 0 0 $X=15402 $Y=5544
XXB19A871F474 GND! VDD! _GENERATED_1432 _GENERATED_1431 278 296 sram_filler $T=15398 4620 0 0 $X=15402 $Y=4620
XXB19A871F475 GND! VDD! _GENERATED_1434 _GENERATED_1433 277 291 sram_filler $T=15398 3696 0 0 $X=15402 $Y=3696
XXB19A871F476 GND! VDD! _GENERATED_1436 _GENERATED_1435 278 296 sram_filler $T=12374 4620 0 0 $X=12378 $Y=4620
XXB19A871F477 GND! VDD! _GENERATED_1438 _GENERATED_1437 277 291 sram_filler $T=12374 3696 0 0 $X=12378 $Y=3696
XXB19A871F478 GND! VDD! _GENERATED_1440 _GENERATED_1439 280 15 sram_filler $T=12374 5544 0 0 $X=12378 $Y=5544
XXB19A871F479 GND! VDD! _GENERATED_1442 _GENERATED_1441 281 15 sram_filler $T=12374 6468 0 0 $X=12378 $Y=6468
XXB19A871F480 GND! VDD! _GENERATED_1444 _GENERATED_1443 277 291 sram_filler $T=9350 3696 0 0 $X=9354 $Y=3696
XXB19A871F481 GND! VDD! _GENERATED_1446 _GENERATED_1445 278 296 sram_filler $T=9350 4620 0 0 $X=9354 $Y=4620
XXB19A871F482 GND! VDD! _GENERATED_1448 _GENERATED_1447 280 15 sram_filler $T=9350 5544 0 0 $X=9354 $Y=5544
XXB19A871F483 GND! VDD! _GENERATED_1450 _GENERATED_1449 281 15 sram_filler $T=9350 6468 0 0 $X=9354 $Y=6468
XXB19A871F484 GND! VDD! GND! _GENERATED_1451 284 300 sram_filler $T=9350 11088 0 0 $X=9354 $Y=11088
XXB19A871F485 GND! VDD! GND! _GENERATED_1452 285 304 sram_filler $T=9350 12012 0 0 $X=9354 $Y=12012
XXB19A871F486 GND! VDD! GND! _GENERATED_1453 287 302 sram_filler $T=9350 13860 0 0 $X=9354 $Y=13860
XXB19A871F487 GND! VDD! GND! _GENERATED_1454 286 303 sram_filler $T=9350 12936 0 0 $X=9354 $Y=12936
XXB19A871F488 GND! VDD! GND! _GENERATED_1455 282 299 sram_filler $T=9350 9240 0 0 $X=9354 $Y=9240
XXB19A871F489 GND! VDD! GND! _GENERATED_1456 283 301 sram_filler $T=9350 10164 0 0 $X=9354 $Y=10164
XXB19A871F490 GND! VDD! GND! _GENERATED_1457 289 297 sram_filler $T=9350 8316 0 0 $X=9354 $Y=8316
XXB19A871F491 GND! VDD! GND! _GENERATED_1458 279 298 sram_filler $T=9350 7392 0 0 $X=9354 $Y=7392
XXB19A871F492 GND! VDD! GND! _GENERATED_1459 284 300 sram_filler $T=12374 11088 0 0 $X=12378 $Y=11088
XXB19A871F493 GND! VDD! GND! _GENERATED_1460 285 304 sram_filler $T=12374 12012 0 0 $X=12378 $Y=12012
XXB19A871F494 GND! VDD! GND! _GENERATED_1461 287 302 sram_filler $T=12374 13860 0 0 $X=12378 $Y=13860
XXB19A871F495 GND! VDD! GND! _GENERATED_1462 286 303 sram_filler $T=12374 12936 0 0 $X=12378 $Y=12936
XXB19A871F496 GND! VDD! GND! _GENERATED_1463 282 299 sram_filler $T=12374 9240 0 0 $X=12378 $Y=9240
XXB19A871F497 GND! VDD! GND! _GENERATED_1464 283 301 sram_filler $T=12374 10164 0 0 $X=12378 $Y=10164
XXB19A871F498 GND! VDD! GND! _GENERATED_1465 289 297 sram_filler $T=12374 8316 0 0 $X=12378 $Y=8316
XXB19A871F499 GND! VDD! GND! _GENERATED_1466 279 298 sram_filler $T=12374 7392 0 0 $X=12378 $Y=7392
XXB19A871F500 GND! VDD! GND! _GENERATED_1467 279 298 sram_filler $T=18422 7392 0 0 $X=18426 $Y=7392
XXB19A871F501 GND! VDD! GND! _GENERATED_1468 289 297 sram_filler $T=18422 8316 0 0 $X=18426 $Y=8316
XXB19A871F502 GND! VDD! GND! _GENERATED_1469 283 301 sram_filler $T=18422 10164 0 0 $X=18426 $Y=10164
XXB19A871F503 GND! VDD! GND! _GENERATED_1470 282 299 sram_filler $T=18422 9240 0 0 $X=18426 $Y=9240
XXB19A871F504 GND! VDD! GND! _GENERATED_1471 286 303 sram_filler $T=18422 12936 0 0 $X=18426 $Y=12936
XXB19A871F505 GND! VDD! GND! _GENERATED_1472 287 302 sram_filler $T=18422 13860 0 0 $X=18426 $Y=13860
XXB19A871F506 GND! VDD! GND! _GENERATED_1473 285 304 sram_filler $T=18422 12012 0 0 $X=18426 $Y=12012
XXB19A871F507 GND! VDD! GND! _GENERATED_1474 284 300 sram_filler $T=18422 11088 0 0 $X=18426 $Y=11088
XXB19A871F508 GND! VDD! GND! _GENERATED_1475 284 300 sram_filler $T=15398 11088 0 0 $X=15402 $Y=11088
XXB19A871F509 GND! VDD! GND! _GENERATED_1476 285 304 sram_filler $T=15398 12012 0 0 $X=15402 $Y=12012
XXB19A871F510 GND! VDD! GND! _GENERATED_1477 287 302 sram_filler $T=15398 13860 0 0 $X=15402 $Y=13860
XXB19A871F511 GND! VDD! GND! _GENERATED_1478 286 303 sram_filler $T=15398 12936 0 0 $X=15402 $Y=12936
XXB19A871F512 GND! VDD! GND! _GENERATED_1479 282 299 sram_filler $T=15398 9240 0 0 $X=15402 $Y=9240
XXB19A871F513 GND! VDD! GND! _GENERATED_1480 283 301 sram_filler $T=15398 10164 0 0 $X=15402 $Y=10164
XXB19A871F514 GND! VDD! GND! _GENERATED_1481 289 297 sram_filler $T=15398 8316 0 0 $X=15402 $Y=8316
XXB19A871F515 GND! VDD! GND! _GENERATED_1482 279 298 sram_filler $T=15398 7392 0 0 $X=15402 $Y=7392
XXB19A871F516 GND! VDD! _GENERATED_1484 _GENERATED_1483 274 293 sram_filler $T=6778 1050 0 180 $X=6330 $Y=460
XXB19A871F517 GND! VDD! _GENERATED_1485 GND! 274 293 sram_filler $T=6442 1050 0 180 $X=5994 $Y=460
XXB19A871F518 GND! VDD! VDD! _GENERATED_1486 274 293 sram_filler $T=6274 1050 0 180 $X=5826 $Y=460
XXB19A871F519 GND! VDD! _GENERATED_1488 _GENERATED_1487 274 293 sram_filler $T=5938 1050 0 180 $X=5489 $Y=460
XXB19A871F520 GND! VDD! _GENERATED_1490 _GENERATED_1489 274 293 sram_filler $T=394 1050 0 180 $X=-53 $Y=460
XXB19A871F521 GND! VDD! _GENERATED_1492 _GENERATED_1491 274 293 sram_filler $T=730 1050 0 180 $X=282 $Y=460
XXB19A871F522 GND! VDD! _GENERATED_1494 _GENERATED_1493 274 293 sram_filler $T=1402 1050 0 180 $X=954 $Y=460
XXB19A871F523 GND! VDD! _GENERATED_1496 _GENERATED_1495 274 293 sram_filler $T=1066 1050 0 180 $X=618 $Y=460
XXB19A871F524 GND! VDD! _GENERATED_1498 _GENERATED_1497 276 294 sram_filler $T=394 1974 0 180 $X=-53 $Y=1384
XXB19A871F525 GND! VDD! _GENERATED_1500 _GENERATED_1499 276 294 sram_filler $T=730 1974 0 180 $X=282 $Y=1384
XXB19A871F526 GND! VDD! _GENERATED_1502 _GENERATED_1501 276 294 sram_filler $T=1402 1974 0 180 $X=954 $Y=1384
XXB19A871F527 GND! VDD! _GENERATED_1504 _GENERATED_1503 276 294 sram_filler $T=1066 1974 0 180 $X=618 $Y=1384
XXB19A871F528 GND! VDD! _GENERATED_1506 _GENERATED_1505 275 295 sram_filler $T=1066 2898 0 180 $X=618 $Y=2308
XXB19A871F529 GND! VDD! _GENERATED_1508 _GENERATED_1507 275 295 sram_filler $T=1402 2898 0 180 $X=954 $Y=2308
XXB19A871F530 GND! VDD! _GENERATED_1510 _GENERATED_1509 275 295 sram_filler $T=730 2898 0 180 $X=282 $Y=2308
XXB19A871F531 GND! VDD! _GENERATED_1512 _GENERATED_1511 275 295 sram_filler $T=394 2898 0 180 $X=-53 $Y=2308
XXB19A871F532 GND! VDD! _GENERATED_1514 _GENERATED_1513 277 292 sram_filler $T=1066 3822 0 180 $X=618 $Y=3232
XXB19A871F533 GND! VDD! _GENERATED_1516 _GENERATED_1515 277 292 sram_filler $T=1402 3822 0 180 $X=954 $Y=3232
XXB19A871F534 GND! VDD! _GENERATED_1518 _GENERATED_1517 277 292 sram_filler $T=730 3822 0 180 $X=282 $Y=3232
XXB19A871F535 GND! VDD! _GENERATED_1520 _GENERATED_1519 277 292 sram_filler $T=394 3822 0 180 $X=-53 $Y=3232
XXB19A871F536 GND! VDD! _GENERATED_1522 _GENERATED_1521 275 295 sram_filler $T=18034 2898 0 180 $X=17586 $Y=2308
XXB19A871F537 GND! VDD! _GENERATED_1524 _GENERATED_1523 275 295 sram_filler $T=18370 2898 0 180 $X=17922 $Y=2308
XXB19A871F538 GND! VDD! 40 _GENERATED_1525 275 295 sram_filler $T=18706 2898 0 180 $X=18258 $Y=2308
XXB19A871F539 GND! VDD! _GENERATED_1527 _GENERATED_1526 275 295 sram_filler $T=16690 2898 0 180 $X=16242 $Y=2308
XXB19A871F540 GND! VDD! _GENERATED_1529 _GENERATED_1528 275 295 sram_filler $T=17026 2898 0 180 $X=16578 $Y=2308
XXB19A871F541 GND! VDD! _GENERATED_1531 _GENERATED_1530 275 295 sram_filler $T=17362 2898 0 180 $X=16914 $Y=2308
XXB19A871F542 GND! VDD! _GENERATED_1533 _GENERATED_1532 275 295 sram_filler $T=17698 2898 0 180 $X=17250 $Y=2308
XXB19A871F543 GND! VDD! VDD! _GENERATED_1534 276 294 sram_filler $T=6610 1974 0 180 $X=6162 $Y=1384
XXB19A871F544 GND! VDD! _GENERATED_1536 _GENERATED_1535 276 294 sram_filler $T=6274 1974 0 180 $X=5826 $Y=1384
XXB19A871F545 GND! VDD! _GENERATED_1538 _GENERATED_1537 276 294 sram_filler $T=5938 1974 0 180 $X=5489 $Y=1384
XXB19A871F546 GND! VDD! _GENERATED_1539 GND! 276 294 sram_filler $T=6778 1974 0 180 $X=6330 $Y=1384
XXB19A871F547 GND! VDD! _GENERATED_1541 _GENERATED_1540 275 295 sram_filler $T=11986 2898 0 180 $X=11538 $Y=2308
XXB19A871F548 GND! VDD! _GENERATED_1543 _GENERATED_1542 275 295 sram_filler $T=12322 2898 0 180 $X=11874 $Y=2308
XXB19A871F549 GND! VDD! _GENERATED_1545 _GENERATED_1544 275 295 sram_filler $T=12658 2898 0 180 $X=12209 $Y=2308
XXB19A871F550 GND! VDD! _GENERATED_1547 _GENERATED_1546 275 295 sram_filler $T=12994 2898 0 180 $X=12546 $Y=2308
XXB19A871F551 GND! VDD! _GENERATED_1549 _GENERATED_1548 275 295 sram_filler $T=13330 2898 0 180 $X=12882 $Y=2308
XXB19A871F552 GND! VDD! _GENERATED_1551 _GENERATED_1550 275 295 sram_filler $T=11314 2898 0 180 $X=10866 $Y=2308
XXB19A871F553 GND! VDD! _GENERATED_1553 _GENERATED_1552 275 295 sram_filler $T=11650 2898 0 180 $X=11202 $Y=2308
XXB19A871F554 GND! VDD! _GENERATED_1555 _GENERATED_1554 275 295 sram_filler $T=13666 2898 0 180 $X=13218 $Y=2308
XXB19A871F555 GND! VDD! _GENERATED_1557 _GENERATED_1556 275 295 sram_filler $T=14002 2898 0 180 $X=13554 $Y=2308
XXB19A871F556 GND! VDD! _GENERATED_1559 _GENERATED_1558 275 295 sram_filler $T=14338 2898 0 180 $X=13890 $Y=2308
XXB19A871F557 GND! VDD! _GENERATED_1561 _GENERATED_1560 275 295 sram_filler $T=14674 2898 0 180 $X=14226 $Y=2308
XXB19A871F558 GND! VDD! _GENERATED_1563 _GENERATED_1562 275 295 sram_filler $T=15010 2898 0 180 $X=14562 $Y=2308
XXB19A871F559 GND! VDD! _GENERATED_1565 _GENERATED_1564 275 295 sram_filler $T=15346 2898 0 180 $X=14898 $Y=2308
XXB19A871F560 GND! VDD! _GENERATED_1567 _GENERATED_1566 275 295 sram_filler $T=16018 2898 0 180 $X=15570 $Y=2308
XXB19A871F561 GND! VDD! _GENERATED_1569 _GENERATED_1568 275 295 sram_filler $T=15682 2898 0 180 $X=15234 $Y=2308
XXB19A871F562 GND! VDD! _GENERATED_1571 _GENERATED_1570 275 295 sram_filler $T=16354 2898 0 180 $X=15905 $Y=2308
XXB19A871F563 GND! VDD! _GENERATED_1573 _GENERATED_1572 275 295 sram_filler $T=9970 2898 0 180 $X=9522 $Y=2308
XXB19A871F564 GND! VDD! _GENERATED_1575 _GENERATED_1574 275 295 sram_filler $T=10306 2898 0 180 $X=9858 $Y=2308
XXB19A871F565 GND! VDD! _GENERATED_1577 _GENERATED_1576 275 295 sram_filler $T=10642 2898 0 180 $X=10193 $Y=2308
XXB19A871F566 GND! VDD! _GENERATED_1579 _GENERATED_1578 275 295 sram_filler $T=10978 2898 0 180 $X=10530 $Y=2308
XXB19A871F567 GND! VDD! _GENERATED_1581 _GENERATED_1580 275 295 sram_filler $T=9634 2898 0 180 $X=9186 $Y=2308
XXB19A871F568 GND! VDD! _GENERATED_1583 _GENERATED_1582 275 295 sram_filler $T=9298 2898 0 180 $X=8850 $Y=2308
XXB19A871F569 GND! VDD! _GENERATED_1585 _GENERATED_1584 275 295 sram_filler $T=8962 2898 0 180 $X=8514 $Y=2308
XXB19A871F570 GND! VDD! _GENERATED_1587 _GENERATED_1586 275 295 sram_filler $T=8626 2898 0 180 $X=8177 $Y=2308
XXB19A871F571 GND! VDD! _GENERATED_1589 _GENERATED_1588 275 295 sram_filler $T=6946 2898 0 180 $X=6497 $Y=2308
XXB19A871F572 GND! VDD! _GENERATED_1591 _GENERATED_1590 275 295 sram_filler $T=6610 2898 0 180 $X=6162 $Y=2308
XXB19A871F573 GND! VDD! _GENERATED_1593 _GENERATED_1592 275 295 sram_filler $T=6274 2898 0 180 $X=5826 $Y=2308
XXB19A871F574 GND! VDD! _GENERATED_1595 _GENERATED_1594 275 295 sram_filler $T=5938 2898 0 180 $X=5489 $Y=2308
XXB19A871F575 GND! VDD! _GENERATED_1597 _GENERATED_1596 275 295 sram_filler $T=8290 2898 0 180 $X=7842 $Y=2308
XXB19A871F576 GND! VDD! _GENERATED_1599 _GENERATED_1598 275 295 sram_filler $T=7954 2898 0 180 $X=7505 $Y=2308
XXB19A871F577 GND! VDD! _GENERATED_1601 _GENERATED_1600 275 295 sram_filler $T=7618 2898 0 180 $X=7170 $Y=2308
XXB19A871F578 GND! VDD! _GENERATED_1603 _GENERATED_1602 275 295 sram_filler $T=7282 2898 0 180 $X=6834 $Y=2308
XXB19A871F579 GND! VDD! _GENERATED_1605 _GENERATED_1604 281 15 sram_filler $T=15850 6594 0 180 $X=15402 $Y=6004
XXB19A871F580 GND! VDD! _GENERATED_1607 _GENERATED_1606 280 296 sram_filler $T=15850 5670 0 180 $X=15402 $Y=5080
XXB19A871F581 GND! VDD! _GENERATED_1609 _GENERATED_1608 278 291 sram_filler $T=15850 4746 0 180 $X=15402 $Y=4156
XXB19A871F582 GND! VDD! _GENERATED_1611 _GENERATED_1610 277 292 sram_filler $T=15850 3822 0 180 $X=15402 $Y=3232
XXB19A871F583 GND! VDD! _GENERATED_1613 _GENERATED_1612 278 291 sram_filler $T=12826 4746 0 180 $X=12378 $Y=4156
XXB19A871F584 GND! VDD! _GENERATED_1615 _GENERATED_1614 277 292 sram_filler $T=12826 3822 0 180 $X=12378 $Y=3232
XXB19A871F585 GND! VDD! _GENERATED_1617 _GENERATED_1616 280 296 sram_filler $T=12826 5670 0 180 $X=12378 $Y=5080
XXB19A871F586 GND! VDD! _GENERATED_1619 _GENERATED_1618 281 15 sram_filler $T=12826 6594 0 180 $X=12378 $Y=6004
XXB19A871F587 GND! VDD! _GENERATED_1621 _GENERATED_1620 277 292 sram_filler $T=9802 3822 0 180 $X=9354 $Y=3232
XXB19A871F588 GND! VDD! _GENERATED_1623 _GENERATED_1622 278 291 sram_filler $T=9802 4746 0 180 $X=9354 $Y=4156
XXB19A871F589 GND! VDD! _GENERATED_1625 _GENERATED_1624 280 296 sram_filler $T=9802 5670 0 180 $X=9354 $Y=5080
XXB19A871F590 GND! VDD! _GENERATED_1627 _GENERATED_1626 281 15 sram_filler $T=9802 6594 0 180 $X=9354 $Y=6004
XXB19A871F591 GND! VDD! VDD! _GENERATED_1628 279 15 sram_filler $T=5938 7518 0 180 $X=5489 $Y=6928
XXB19A871F592 GND! VDD! _GENERATED_1629 GND! 279 15 sram_filler $T=6106 7518 0 180 $X=5657 $Y=6928
XXB19A871F593 GND! VDD! _GENERATED_1631 _GENERATED_1630 279 15 sram_filler $T=6442 7518 0 180 $X=5994 $Y=6928
XXB19A871F594 GND! VDD! VDD! _GENERATED_1632 278 291 sram_filler $T=394 4746 0 180 $X=-53 $Y=4156
XXB19A871F595 GND! VDD! _GENERATED_1634 _GENERATED_1633 278 291 sram_filler $T=2914 4746 0 180 $X=2466 $Y=4156
XXB19A871F596 GND! VDD! _GENERATED_1636 _GENERATED_1635 278 291 sram_filler $T=2578 4746 0 180 $X=2130 $Y=4156
XXB19A871F597 GND! VDD! _GENERATED_1638 _GENERATED_1637 278 291 sram_filler $T=1906 4746 0 180 $X=1458 $Y=4156
XXB19A871F598 GND! VDD! _GENERATED_1640 _GENERATED_1639 278 291 sram_filler $T=2242 4746 0 180 $X=1794 $Y=4156
XXB19A871F599 GND! VDD! _GENERATED_1642 _GENERATED_1641 278 291 sram_filler $T=1234 4746 0 180 $X=786 $Y=4156
XXB19A871F600 GND! VDD! _GENERATED_1644 _GENERATED_1643 278 291 sram_filler $T=1570 4746 0 180 $X=1122 $Y=4156
XXB19A871F601 GND! VDD! _GENERATED_1645 GND! 278 291 sram_filler $T=562 4746 0 180 $X=114 $Y=4156
XXB19A871F602 GND! VDD! _GENERATED_1647 _GENERATED_1646 278 291 sram_filler $T=898 4746 0 180 $X=450 $Y=4156
XXB19A871F603 GND! VDD! _GENERATED_1649 _GENERATED_1648 278 291 sram_filler $T=3586 4746 0 180 $X=3138 $Y=4156
XXB19A871F604 GND! VDD! _GENERATED_1651 _GENERATED_1650 278 291 sram_filler $T=3250 4746 0 180 $X=2802 $Y=4156
XXB19A871F605 GND! VDD! _GENERATED_1653 _GENERATED_1652 278 291 sram_filler $T=4258 4746 0 180 $X=3810 $Y=4156
XXB19A871F606 GND! VDD! _GENERATED_1655 _GENERATED_1654 278 291 sram_filler $T=3922 4746 0 180 $X=3474 $Y=4156
XXB19A871F607 GND! VDD! _GENERATED_1657 _GENERATED_1656 278 291 sram_filler $T=4930 4746 0 180 $X=4481 $Y=4156
XXB19A871F608 GND! VDD! _GENERATED_1659 _GENERATED_1658 278 291 sram_filler $T=4594 4746 0 180 $X=4146 $Y=4156
XXB19A871F609 GND! VDD! _GENERATED_1661 _GENERATED_1660 278 291 sram_filler $T=5266 4746 0 180 $X=4818 $Y=4156
XXB19A871F610 GND! VDD! _GENERATED_1663 _GENERATED_1662 278 291 sram_filler $T=5602 4746 0 180 $X=5154 $Y=4156
XXB19A871F611 GND! VDD! _GENERATED_1665 _GENERATED_1664 279 15 sram_filler $T=6778 7518 0 180 $X=6330 $Y=6928
XXB19A871F612 GND! VDD! GND! _GENERATED_1666 285 300 sram_filler $T=9350 12138 1 0 $X=9354 $Y=11548
XXB19A871F613 GND! VDD! GND! _GENERATED_1667 286 304 sram_filler $T=9350 13062 1 0 $X=9354 $Y=12472
XXB19A871F614 GND! VDD! GND! _GENERATED_1668 288 302 sram_filler $T=9350 14910 1 0 $X=9354 $Y=14320
XXB19A871F615 GND! VDD! GND! _GENERATED_1669 287 303 sram_filler $T=9350 13986 1 0 $X=9354 $Y=13396
XXB19A871F616 GND! VDD! GND! _GENERATED_1670 283 299 sram_filler $T=9350 10290 1 0 $X=9354 $Y=9700
XXB19A871F617 GND! VDD! GND! _GENERATED_1671 284 301 sram_filler $T=9350 11214 1 0 $X=9354 $Y=10624
XXB19A871F618 GND! VDD! GND! _GENERATED_1672 282 297 sram_filler $T=9350 9366 1 0 $X=9354 $Y=8776
XXB19A871F619 GND! VDD! GND! _GENERATED_1673 289 298 sram_filler $T=9350 8442 1 0 $X=9354 $Y=7852
XXB19A871F620 GND! VDD! GND! _GENERATED_1674 285 300 sram_filler $T=12374 12138 1 0 $X=12378 $Y=11548
XXB19A871F621 GND! VDD! GND! _GENERATED_1675 286 304 sram_filler $T=12374 13062 1 0 $X=12378 $Y=12472
XXB19A871F622 GND! VDD! GND! _GENERATED_1676 288 302 sram_filler $T=12374 14910 1 0 $X=12378 $Y=14320
XXB19A871F623 GND! VDD! GND! _GENERATED_1677 287 303 sram_filler $T=12374 13986 1 0 $X=12378 $Y=13396
XXB19A871F624 GND! VDD! GND! _GENERATED_1678 283 299 sram_filler $T=12374 10290 1 0 $X=12378 $Y=9700
XXB19A871F625 GND! VDD! GND! _GENERATED_1679 284 301 sram_filler $T=12374 11214 1 0 $X=12378 $Y=10624
XXB19A871F626 GND! VDD! GND! _GENERATED_1680 282 297 sram_filler $T=12374 9366 1 0 $X=12378 $Y=8776
XXB19A871F627 GND! VDD! GND! _GENERATED_1681 289 298 sram_filler $T=12374 8442 1 0 $X=12378 $Y=7852
XXB19A871F628 GND! VDD! GND! _GENERATED_1682 289 298 sram_filler $T=18422 8442 1 0 $X=18426 $Y=7852
XXB19A871F629 GND! VDD! GND! _GENERATED_1683 282 297 sram_filler $T=18422 9366 1 0 $X=18426 $Y=8776
XXB19A871F630 GND! VDD! GND! _GENERATED_1684 284 301 sram_filler $T=18422 11214 1 0 $X=18426 $Y=10624
XXB19A871F631 GND! VDD! GND! _GENERATED_1685 283 299 sram_filler $T=18422 10290 1 0 $X=18426 $Y=9700
XXB19A871F632 GND! VDD! GND! _GENERATED_1686 287 303 sram_filler $T=18422 13986 1 0 $X=18426 $Y=13396
XXB19A871F633 GND! VDD! GND! _GENERATED_1687 288 302 sram_filler $T=18422 14910 1 0 $X=18426 $Y=14320
XXB19A871F634 GND! VDD! GND! _GENERATED_1688 286 304 sram_filler $T=18422 13062 1 0 $X=18426 $Y=12472
XXB19A871F635 GND! VDD! GND! _GENERATED_1689 285 300 sram_filler $T=18422 12138 1 0 $X=18426 $Y=11548
XXB19A871F636 GND! VDD! GND! _GENERATED_1690 285 300 sram_filler $T=15398 12138 1 0 $X=15402 $Y=11548
XXB19A871F637 GND! VDD! GND! _GENERATED_1691 286 304 sram_filler $T=15398 13062 1 0 $X=15402 $Y=12472
XXB19A871F638 GND! VDD! GND! _GENERATED_1692 288 302 sram_filler $T=15398 14910 1 0 $X=15402 $Y=14320
XXB19A871F639 GND! VDD! GND! _GENERATED_1693 287 303 sram_filler $T=15398 13986 1 0 $X=15402 $Y=13396
XXB19A871F640 GND! VDD! GND! _GENERATED_1694 283 299 sram_filler $T=15398 10290 1 0 $X=15402 $Y=9700
XXB19A871F641 GND! VDD! GND! _GENERATED_1695 284 301 sram_filler $T=15398 11214 1 0 $X=15402 $Y=10624
XXB19A871F642 GND! VDD! GND! _GENERATED_1696 282 297 sram_filler $T=15398 9366 1 0 $X=15402 $Y=8776
XXB19A871F643 GND! VDD! GND! _GENERATED_1697 289 298 sram_filler $T=15398 8442 1 0 $X=15402 $Y=7852
XXB19A871F644 GND! VDD! GND! 15 379 157 14 119 194 120 282 
+	283 299 sram_6t $T=6690 9240 0 0 $X=6666 $Y=9240
XXB19A871F645 GND! VDD! GND! 9 347 493 8 115 150 116 279 
+	289 298 sram_6t $T=8706 7392 0 0 $X=8682 $Y=7392
XXB19A871F646 GND! VDD! GND! 11 348 494 10 115 151 116 279 
+	289 298 sram_6t $T=8034 7392 0 0 $X=8010 $Y=7392
XXB19A871F647 GND! VDD! GND! 13 349 495 12 115 152 116 279 
+	289 298 sram_6t $T=7362 7392 0 0 $X=7338 $Y=7392
XXB19A871F648 GND! VDD! GND! 13 350 152 12 116 153 119 289 
+	282 297 sram_6t $T=7362 8316 0 0 $X=7338 $Y=8316
XXB19A871F649 GND! VDD! GND! 11 351 151 10 116 154 119 289 
+	282 297 sram_6t $T=8034 8316 0 0 $X=8010 $Y=8316
XXB19A871F650 GND! VDD! GND! 9 352 150 8 116 155 119 289 
+	282 297 sram_6t $T=8706 8316 0 0 $X=8682 $Y=8316
XXB19A871F651 GND! VDD! GND! 15 353 496 14 115 156 116 279 
+	289 298 sram_6t $T=6690 7392 0 0 $X=6666 $Y=7392
XXB19A871F652 GND! VDD! GND! 15 354 156 14 116 157 119 289 
+	282 297 sram_6t $T=6690 8316 0 0 $X=6666 $Y=8316
XXB19A871F653 GND! VDD! GND! 13 380 153 12 119 195 120 282 
+	283 299 sram_6t $T=7362 9240 0 0 $X=7338 $Y=9240
XXB19A871F654 GND! VDD! GND! 11 381 154 10 119 196 120 282 
+	283 299 sram_6t $T=8034 9240 0 0 $X=8010 $Y=9240
XXB19A871F655 GND! VDD! GND! 9 382 155 8 119 197 120 282 
+	283 299 sram_6t $T=8706 9240 0 0 $X=8682 $Y=9240
XXB19A871F656 GND! VDD! GND! 15 383 194 14 120 198 121 283 
+	284 301 sram_6t $T=6690 10164 0 0 $X=6666 $Y=10164
XXB19A871F657 GND! VDD! GND! 9 384 197 8 120 199 121 283 
+	284 301 sram_6t $T=8706 10164 0 0 $X=8682 $Y=10164
XXB19A871F658 GND! VDD! GND! 11 385 196 10 120 200 121 283 
+	284 301 sram_6t $T=8034 10164 0 0 $X=8010 $Y=10164
XXB19A871F659 GND! VDD! GND! 13 386 195 12 120 201 121 283 
+	284 301 sram_6t $T=7362 10164 0 0 $X=7338 $Y=10164
XXB19A871F660 GND! VDD! GND! 9 387 199 8 121 202 122 284 
+	285 300 sram_6t $T=8706 11088 0 0 $X=8682 $Y=11088
XXB19A871F661 GND! VDD! GND! 11 388 200 10 121 203 122 284 
+	285 300 sram_6t $T=8034 11088 0 0 $X=8010 $Y=11088
XXB19A871F662 GND! VDD! GND! 13 389 201 12 121 204 122 284 
+	285 300 sram_6t $T=7362 11088 0 0 $X=7338 $Y=11088
XXB19A871F663 GND! VDD! GND! 15 390 198 14 121 205 122 284 
+	285 300 sram_6t $T=6690 11088 0 0 $X=6666 $Y=11088
XXB19A871F664 GND! VDD! GND! 13 427 204 12 122 206 123 285 
+	286 304 sram_6t $T=7362 12012 0 0 $X=7338 $Y=12012
XXB19A871F665 GND! VDD! GND! 11 428 203 10 122 207 123 285 
+	286 304 sram_6t $T=8034 12012 0 0 $X=8010 $Y=12012
XXB19A871F666 GND! VDD! GND! 9 429 202 8 122 208 123 285 
+	286 304 sram_6t $T=8706 12012 0 0 $X=8682 $Y=12012
XXB19A871F667 GND! VDD! GND! 15 430 205 14 122 209 123 285 
+	286 304 sram_6t $T=6690 12012 0 0 $X=6666 $Y=12012
XXB19A871F668 GND! VDD! GND! 15 431 209 14 123 210 124 286 
+	287 303 sram_6t $T=6690 12936 0 0 $X=6666 $Y=12936
XXB19A871F669 GND! VDD! GND! 13 432 206 12 123 211 124 286 
+	287 303 sram_6t $T=7362 12936 0 0 $X=7338 $Y=12936
XXB19A871F670 GND! VDD! GND! 11 433 207 10 123 212 124 286 
+	287 303 sram_6t $T=8034 12936 0 0 $X=8010 $Y=12936
XXB19A871F671 GND! VDD! GND! 9 434 208 8 123 213 124 286 
+	287 303 sram_6t $T=8706 12936 0 0 $X=8682 $Y=12936
XXB19A871F672 GND! VDD! GND! 15 435 210 14 124 518 519 287 
+	288 302 sram_6t $T=6690 13860 0 0 $X=6666 $Y=13860
XXB19A871F673 GND! VDD! GND! 9 436 213 8 124 524 525 287 
+	288 302 sram_6t $T=8706 13860 0 0 $X=8682 $Y=13860
XXB19A871F674 GND! VDD! GND! 11 437 212 10 124 522 523 287 
+	288 302 sram_6t $T=8034 13860 0 0 $X=8010 $Y=13860
XXB19A871F675 GND! VDD! GND! 13 438 211 12 124 520 521 287 
+	288 302 sram_6t $T=7362 13860 0 0 $X=7338 $Y=13860
XXB19A871F676 GND! VDD! GND! 18 439 214 19 124 528 529 287 
+	288 302 sram_6t $T=10386 13860 0 0 $X=10362 $Y=13860
XXB19A871F677 GND! VDD! GND! 20 440 215 21 124 530 531 287 
+	288 302 sram_6t $T=11058 13860 0 0 $X=11034 $Y=13860
XXB19A871F678 GND! VDD! GND! 22 441 216 23 124 532 533 287 
+	288 302 sram_6t $T=11730 13860 0 0 $X=11706 $Y=13860
XXB19A871F679 GND! VDD! GND! 17 442 217 16 124 526 527 287 
+	288 302 sram_6t $T=9714 13860 0 0 $X=9690 $Y=13860
XXB19A871F680 GND! VDD! GND! 22 443 218 23 123 216 124 286 
+	287 303 sram_6t $T=11730 12936 0 0 $X=11706 $Y=12936
XXB19A871F681 GND! VDD! GND! 20 444 219 21 123 215 124 286 
+	287 303 sram_6t $T=11058 12936 0 0 $X=11034 $Y=12936
XXB19A871F682 GND! VDD! GND! 18 445 220 19 123 214 124 286 
+	287 303 sram_6t $T=10386 12936 0 0 $X=10362 $Y=12936
XXB19A871F683 GND! VDD! GND! 17 446 221 16 123 217 124 286 
+	287 303 sram_6t $T=9714 12936 0 0 $X=9690 $Y=12936
XXB19A871F684 GND! VDD! GND! 17 447 222 16 122 221 123 285 
+	286 304 sram_6t $T=9714 12012 0 0 $X=9690 $Y=12012
XXB19A871F685 GND! VDD! GND! 22 448 223 23 122 218 123 285 
+	286 304 sram_6t $T=11730 12012 0 0 $X=11706 $Y=12012
XXB19A871F686 GND! VDD! GND! 20 449 224 21 122 219 123 285 
+	286 304 sram_6t $T=11058 12012 0 0 $X=11034 $Y=12012
XXB19A871F687 GND! VDD! GND! 18 450 225 19 122 220 123 285 
+	286 304 sram_6t $T=10386 12012 0 0 $X=10362 $Y=12012
XXB19A871F688 GND! VDD! GND! 17 391 226 16 121 222 122 284 
+	285 300 sram_6t $T=9714 11088 0 0 $X=9690 $Y=11088
XXB19A871F689 GND! VDD! GND! 18 392 227 19 121 225 122 284 
+	285 300 sram_6t $T=10386 11088 0 0 $X=10362 $Y=11088
XXB19A871F690 GND! VDD! GND! 20 393 228 21 121 224 122 284 
+	285 300 sram_6t $T=11058 11088 0 0 $X=11034 $Y=11088
XXB19A871F691 GND! VDD! GND! 22 394 229 23 121 223 122 284 
+	285 300 sram_6t $T=11730 11088 0 0 $X=11706 $Y=11088
XXB19A871F692 GND! VDD! GND! 18 395 230 19 120 227 121 283 
+	284 301 sram_6t $T=10386 10164 0 0 $X=10362 $Y=10164
XXB19A871F693 GND! VDD! GND! 20 396 231 21 120 228 121 283 
+	284 301 sram_6t $T=11058 10164 0 0 $X=11034 $Y=10164
XXB19A871F694 GND! VDD! GND! 22 397 232 23 120 229 121 283 
+	284 301 sram_6t $T=11730 10164 0 0 $X=11706 $Y=10164
XXB19A871F695 GND! VDD! GND! 17 398 233 16 120 226 121 283 
+	284 301 sram_6t $T=9714 10164 0 0 $X=9690 $Y=10164
XXB19A871F696 GND! VDD! GND! 22 399 169 23 119 232 120 282 
+	283 299 sram_6t $T=11730 9240 0 0 $X=11706 $Y=9240
XXB19A871F697 GND! VDD! GND! 20 400 167 21 119 231 120 282 
+	283 299 sram_6t $T=11058 9240 0 0 $X=11034 $Y=9240
XXB19A871F698 GND! VDD! GND! 18 401 165 19 119 230 120 282 
+	283 299 sram_6t $T=10386 9240 0 0 $X=10362 $Y=9240
XXB19A871F699 GND! VDD! GND! 17 402 163 16 119 233 120 282 
+	283 299 sram_6t $T=9714 9240 0 0 $X=9690 $Y=9240
XXB19A871F700 GND! VDD! GND! 17 355 162 16 116 163 119 289 
+	282 297 sram_6t $T=9714 8316 0 0 $X=9690 $Y=8316
XXB19A871F701 GND! VDD! GND! 18 356 164 19 116 165 119 289 
+	282 297 sram_6t $T=10386 8316 0 0 $X=10362 $Y=8316
XXB19A871F702 GND! VDD! GND! 20 357 166 21 116 167 119 289 
+	282 297 sram_6t $T=11058 8316 0 0 $X=11034 $Y=8316
XXB19A871F703 GND! VDD! GND! 22 358 168 23 116 169 119 289 
+	282 297 sram_6t $T=11730 8316 0 0 $X=11706 $Y=8316
XXB19A871F704 GND! VDD! GND! 22 359 497 23 115 168 116 279 
+	289 298 sram_6t $T=11730 7392 0 0 $X=11706 $Y=7392
XXB19A871F705 GND! VDD! GND! 20 360 498 21 115 166 116 279 
+	289 298 sram_6t $T=11058 7392 0 0 $X=11034 $Y=7392
XXB19A871F706 GND! VDD! GND! 18 361 499 19 115 164 116 279 
+	289 298 sram_6t $T=10386 7392 0 0 $X=10362 $Y=7392
XXB19A871F707 GND! VDD! GND! 17 362 500 16 115 162 116 279 
+	289 298 sram_6t $T=9714 7392 0 0 $X=9690 $Y=7392
XXB19A871F708 GND! VDD! GND! 39 363 186 38 116 187 119 289 
+	282 297 sram_6t $T=17778 8316 0 0 $X=17753 $Y=8316
XXB19A871F709 GND! VDD! GND! 37 364 188 36 116 189 119 289 
+	282 297 sram_6t $T=17106 8316 0 0 $X=17082 $Y=8316
XXB19A871F710 GND! VDD! GND! 35 365 190 34 116 191 119 289 
+	282 297 sram_6t $T=16434 8316 0 0 $X=16410 $Y=8316
XXB19A871F711 GND! VDD! GND! 33 366 192 32 116 193 119 289 
+	282 297 sram_6t $T=15762 8316 0 0 $X=15738 $Y=8316
XXB19A871F712 GND! VDD! GND! 33 403 193 32 119 254 120 282 
+	283 299 sram_6t $T=15762 9240 0 0 $X=15738 $Y=9240
XXB19A871F713 GND! VDD! GND! 35 404 191 34 119 255 120 282 
+	283 299 sram_6t $T=16434 9240 0 0 $X=16410 $Y=9240
XXB19A871F714 GND! VDD! GND! 37 405 189 36 119 256 120 282 
+	283 299 sram_6t $T=17106 9240 0 0 $X=17082 $Y=9240
XXB19A871F715 GND! VDD! GND! 39 406 187 38 119 257 120 282 
+	283 299 sram_6t $T=17778 9240 0 0 $X=17753 $Y=9240
XXB19A871F716 GND! VDD! GND! 33 407 254 32 120 258 121 283 
+	284 301 sram_6t $T=15762 10164 0 0 $X=15738 $Y=10164
XXB19A871F717 GND! VDD! GND! 39 408 257 38 120 259 121 283 
+	284 301 sram_6t $T=17778 10164 0 0 $X=17753 $Y=10164
XXB19A871F718 GND! VDD! GND! 37 409 256 36 120 260 121 283 
+	284 301 sram_6t $T=17106 10164 0 0 $X=17082 $Y=10164
XXB19A871F719 GND! VDD! GND! 35 410 255 34 120 261 121 283 
+	284 301 sram_6t $T=16434 10164 0 0 $X=16410 $Y=10164
XXB19A871F720 GND! VDD! GND! 39 411 259 38 121 262 122 284 
+	285 300 sram_6t $T=17778 11088 0 0 $X=17753 $Y=11088
XXB19A871F721 GND! VDD! GND! 37 412 260 36 121 263 122 284 
+	285 300 sram_6t $T=17106 11088 0 0 $X=17082 $Y=11088
XXB19A871F722 GND! VDD! GND! 35 413 261 34 121 264 122 284 
+	285 300 sram_6t $T=16434 11088 0 0 $X=16410 $Y=11088
XXB19A871F723 GND! VDD! GND! 33 414 258 32 121 265 122 284 
+	285 300 sram_6t $T=15762 11088 0 0 $X=15738 $Y=11088
XXB19A871F724 GND! VDD! GND! 35 451 264 34 122 266 123 285 
+	286 304 sram_6t $T=16434 12012 0 0 $X=16410 $Y=12012
XXB19A871F725 GND! VDD! GND! 37 452 263 36 122 267 123 285 
+	286 304 sram_6t $T=17106 12012 0 0 $X=17082 $Y=12012
XXB19A871F726 GND! VDD! GND! 39 453 262 38 122 268 123 285 
+	286 304 sram_6t $T=17778 12012 0 0 $X=17753 $Y=12012
XXB19A871F727 GND! VDD! GND! 33 454 265 32 122 269 123 285 
+	286 304 sram_6t $T=15762 12012 0 0 $X=15738 $Y=12012
XXB19A871F728 GND! VDD! GND! 33 455 269 32 123 270 124 286 
+	287 303 sram_6t $T=15762 12936 0 0 $X=15738 $Y=12936
XXB19A871F729 GND! VDD! GND! 35 456 266 34 123 271 124 286 
+	287 303 sram_6t $T=16434 12936 0 0 $X=16410 $Y=12936
XXB19A871F730 GND! VDD! GND! 37 457 267 36 123 272 124 286 
+	287 303 sram_6t $T=17106 12936 0 0 $X=17082 $Y=12936
XXB19A871F731 GND! VDD! GND! 39 458 268 38 123 273 124 286 
+	287 303 sram_6t $T=17778 12936 0 0 $X=17753 $Y=12936
XXB19A871F732 GND! VDD! GND! 33 459 270 32 124 542 543 287 
+	288 302 sram_6t $T=15762 13860 0 0 $X=15738 $Y=13860
XXB19A871F733 GND! VDD! GND! 39 460 273 38 124 548 549 287 
+	288 302 sram_6t $T=17778 13860 0 0 $X=17753 $Y=13860
XXB19A871F734 GND! VDD! GND! 37 461 272 36 124 546 547 287 
+	288 302 sram_6t $T=17106 13860 0 0 $X=17082 $Y=13860
XXB19A871F735 GND! VDD! GND! 35 462 271 34 124 544 545 287 
+	288 302 sram_6t $T=16434 13860 0 0 $X=16410 $Y=13860
XXB19A871F736 GND! VDD! GND! 30 463 234 31 124 540 541 287 
+	288 302 sram_6t $T=14754 13860 0 0 $X=14730 $Y=13860
XXB19A871F737 GND! VDD! GND! 30 464 235 31 123 234 124 286 
+	287 303 sram_6t $T=14754 12936 0 0 $X=14730 $Y=12936
XXB19A871F738 GND! VDD! GND! 30 465 236 31 122 235 123 285 
+	286 304 sram_6t $T=14754 12012 0 0 $X=14730 $Y=12012
XXB19A871F739 GND! VDD! GND! 30 415 237 31 121 236 122 284 
+	285 300 sram_6t $T=14754 11088 0 0 $X=14730 $Y=11088
XXB19A871F740 GND! VDD! GND! 30 416 238 31 120 237 121 283 
+	284 301 sram_6t $T=14754 10164 0 0 $X=14730 $Y=10164
XXB19A871F741 GND! VDD! GND! 30 417 175 31 119 238 120 282 
+	283 299 sram_6t $T=14754 9240 0 0 $X=14730 $Y=9240
XXB19A871F742 GND! VDD! GND! 30 367 174 31 116 175 119 289 
+	282 297 sram_6t $T=14754 8316 0 0 $X=14730 $Y=8316
XXB19A871F743 GND! VDD! GND! 33 368 503 32 115 192 116 279 
+	289 298 sram_6t $T=15762 7392 0 0 $X=15738 $Y=7392
XXB19A871F744 GND! VDD! GND! 35 369 504 34 115 190 116 279 
+	289 298 sram_6t $T=16434 7392 0 0 $X=16410 $Y=7392
XXB19A871F745 GND! VDD! GND! 37 370 505 36 115 188 116 279 
+	289 298 sram_6t $T=17106 7392 0 0 $X=17082 $Y=7392
XXB19A871F746 GND! VDD! GND! 39 371 506 38 115 186 116 279 
+	289 298 sram_6t $T=17778 7392 0 0 $X=17753 $Y=7392
XXB19A871F747 GND! VDD! GND! 27 466 239 26 124 536 537 287 
+	288 302 sram_6t $T=13410 13860 0 0 $X=13386 $Y=13860
XXB19A871F748 GND! VDD! GND! 25 467 240 24 124 538 539 287 
+	288 302 sram_6t $T=14082 13860 0 0 $X=14058 $Y=13860
XXB19A871F749 GND! VDD! GND! 29 468 241 28 124 534 535 287 
+	288 302 sram_6t $T=12738 13860 0 0 $X=12714 $Y=13860
XXB19A871F750 GND! VDD! GND! 25 469 242 24 123 240 124 286 
+	287 303 sram_6t $T=14082 12936 0 0 $X=14058 $Y=12936
XXB19A871F751 GND! VDD! GND! 27 470 243 26 123 239 124 286 
+	287 303 sram_6t $T=13410 12936 0 0 $X=13386 $Y=12936
XXB19A871F752 GND! VDD! GND! 29 471 244 28 123 241 124 286 
+	287 303 sram_6t $T=12738 12936 0 0 $X=12714 $Y=12936
XXB19A871F753 GND! VDD! GND! 29 472 245 28 122 244 123 285 
+	286 304 sram_6t $T=12738 12012 0 0 $X=12714 $Y=12012
XXB19A871F754 GND! VDD! GND! 25 473 246 24 122 242 123 285 
+	286 304 sram_6t $T=14082 12012 0 0 $X=14058 $Y=12012
XXB19A871F755 GND! VDD! GND! 27 474 247 26 122 243 123 285 
+	286 304 sram_6t $T=13410 12012 0 0 $X=13386 $Y=12012
XXB19A871F756 GND! VDD! GND! 29 418 248 28 121 245 122 284 
+	285 300 sram_6t $T=12738 11088 0 0 $X=12714 $Y=11088
XXB19A871F757 GND! VDD! GND! 27 419 249 26 121 247 122 284 
+	285 300 sram_6t $T=13410 11088 0 0 $X=13386 $Y=11088
XXB19A871F758 GND! VDD! GND! 25 420 250 24 121 246 122 284 
+	285 300 sram_6t $T=14082 11088 0 0 $X=14058 $Y=11088
XXB19A871F759 GND! VDD! GND! 27 421 251 26 120 249 121 283 
+	284 301 sram_6t $T=13410 10164 0 0 $X=13386 $Y=10164
XXB19A871F760 GND! VDD! GND! 25 422 252 24 120 250 121 283 
+	284 301 sram_6t $T=14082 10164 0 0 $X=14058 $Y=10164
XXB19A871F761 GND! VDD! GND! 29 423 253 28 120 248 121 283 
+	284 301 sram_6t $T=12738 10164 0 0 $X=12714 $Y=10164
XXB19A871F762 GND! VDD! GND! 25 424 181 24 119 252 120 282 
+	283 299 sram_6t $T=14082 9240 0 0 $X=14058 $Y=9240
XXB19A871F763 GND! VDD! GND! 27 425 179 26 119 251 120 282 
+	283 299 sram_6t $T=13410 9240 0 0 $X=13386 $Y=9240
XXB19A871F764 GND! VDD! GND! 29 426 177 28 119 253 120 282 
+	283 299 sram_6t $T=12738 9240 0 0 $X=12714 $Y=9240
XXB19A871F765 GND! VDD! GND! 29 372 176 28 116 177 119 289 
+	282 297 sram_6t $T=12738 8316 0 0 $X=12714 $Y=8316
XXB19A871F766 GND! VDD! GND! 27 373 178 26 116 179 119 289 
+	282 297 sram_6t $T=13410 8316 0 0 $X=13386 $Y=8316
XXB19A871F767 GND! VDD! GND! 25 374 180 24 116 181 119 289 
+	282 297 sram_6t $T=14082 8316 0 0 $X=14058 $Y=8316
XXB19A871F768 GND! VDD! GND! 30 375 507 31 115 174 116 279 
+	289 298 sram_6t $T=14754 7392 0 0 $X=14730 $Y=7392
XXB19A871F769 GND! VDD! GND! 25 376 508 24 115 180 116 279 
+	289 298 sram_6t $T=14082 7392 0 0 $X=14058 $Y=7392
XXB19A871F770 GND! VDD! GND! 27 377 501 26 115 178 116 279 
+	289 298 sram_6t $T=13410 7392 0 0 $X=13386 $Y=7392
XXB19A871F771 GND! VDD! GND! 29 378 502 28 115 176 116 279 
+	289 298 sram_6t $T=12738 7392 0 0 $X=12714 $Y=7392
.ends memory_array_static_column_decoder_test
