* PEX netlist file	Wed Apr 16 22:21:51 2025	agen_unit
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 2
.subckt inv 2 3 4 5 7 8
*.floating_nets 6
.ends inv
.subckt nand 2 3 4 5 6 7 8 9 12 13
*.floating_nets 10 11
.ends nand
.subckt sram_filler 2 3 4 5 6 7
.ends sram_filler
.subckt nor 2 3 4 5 6 7 8 9 10 11 12
.ends nor
.subckt invx4 2 3 4 5 6 7 8 9 10 11 12
+	13
.ends invx4

* Hierarchy Level 1
.subckt Demux 2 3 4 5 6 7 8 9 10 11 12
+	13 14 16
MM1 10 8 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1398 $Y=315  $PIN_XY=1428,378,1398,315,1368,378 $DEVICE_ID=1001
MM2 8 5 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=894 $Y=315  $PIN_XY=924,378,894,315,864,378 $DEVICE_ID=1001
MM3 15 7 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=726 $Y=315  $PIN_XY=756,378,726,315,696,378 $DEVICE_ID=1001
XXCE9F2C6675 2 3 6 5 12 13 inv $T=0 462 0 0 $X=0 $Y=462
XXCE9F2C6676 2 3 11 9 12 13 inv $T=1176 462 0 0 $X=1176 $Y=462
XXCE9F2C6677 2 4 10 8 12 14 inv $T=1176 588 1 0 $X=1176 $Y=-2
XXCE9F2C6678 2 4 _GENERATED_17 2 12 14 sram_filler $T=616 588 0 180 $X=167 $Y=-2
XXCE9F2C6679 2 4 4 _GENERATED_18 12 14 sram_filler $T=448 588 0 180 $X=0 $Y=-2
XXCE9F2C6680 2 3 9 7 6 7 5 16 12 13 nand $T=86 234 0 0 $X=504 $Y=462
XXCE9F2C6681 2 4 8 7 5 7 6 15 12 14 nand $T=86 816 1 0 $X=504 $Y=-2
.ends Demux

* Hierarchy Level 0

* Top of hierarchy  cell=agen_unit
.subckt agen_unit GND! VDD! 4 5 6 7 8 9 10 11 WEN
+	13 14 15 16 17 18 WS0 RS1 RS1BAR WS1 WS1BAR
+	RS0 RS0BAR WS0BAR 27 28 29 A1 A0
*.floating_nets 57 58 59 60 61 62 63 64 65 66 67
*+	_GENERATED_918 _GENERATED_919
MM1 GND! 16 WS0BAR nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=1916  $PIN_XY=3782,1832,3752,1916,3722,1832 $DEVICE_ID=1001
MM2 GND! 18 WS0 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=1454  $PIN_XY=3782,1538,3752,1454,3722,1538 $DEVICE_ID=1001
MM3 GND! 14 RS0BAR nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=992  $PIN_XY=3782,908,3752,992,3722,908 $DEVICE_ID=1001
MM4 GND! 27 RS0 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=530  $PIN_XY=3782,614,3752,530,3722,614 $DEVICE_ID=1001
MM5 GND! 17 WS1BAR nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=68  $PIN_XY=3782,-16,3752,68,3722,-16 $DEVICE_ID=1001
MM6 GND! 15 WS1 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=-394  $PIN_XY=3782,-310,3752,-394,3722,-310 $DEVICE_ID=1001
MM7 GND! 29 RS1BAR nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=-856  $PIN_XY=3782,-940,3752,-856,3722,-940 $DEVICE_ID=1001
MM8 GND! 28 RS1 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3752 $Y=-1318  $PIN_XY=3782,-1234,3752,-1318,3722,-1234 $DEVICE_ID=1001
MM9 WS0BAR 16 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=1916  $PIN_XY=3614,1832,3584,1916,3554,1832 $DEVICE_ID=1001
MM10 WS0 18 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=1454  $PIN_XY=3614,1538,3584,1454,3554,1538 $DEVICE_ID=1001
MM11 RS0BAR 14 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=992  $PIN_XY=3614,908,3584,992,3554,908 $DEVICE_ID=1001
MM12 RS0 27 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=530  $PIN_XY=3614,614,3584,530,3554,614 $DEVICE_ID=1001
MM13 WS1BAR 17 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=68  $PIN_XY=3614,-16,3584,68,3554,-16 $DEVICE_ID=1001
MM14 WS1 15 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-394  $PIN_XY=3614,-310,3584,-394,3554,-310 $DEVICE_ID=1001
MM15 RS1BAR 29 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-856  $PIN_XY=3614,-940,3584,-856,3554,-940 $DEVICE_ID=1001
MM16 RS1 28 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-1318  $PIN_XY=3614,-1234,3584,-1318,3554,-1234 $DEVICE_ID=1001
MM17 GND! 5 14 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=971  $PIN_XY=3278,908,3248,971,3218,908 $DEVICE_ID=1001
MM18 GND! 10 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=551  $PIN_XY=3278,614,3248,551,3218,614 $DEVICE_ID=1001
MM19 GND! 4 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=-877  $PIN_XY=3278,-940,3248,-877,3218,-940 $DEVICE_ID=1001
MM20 GND! 8 28 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=-1318  $PIN_XY=3278,-1234,3248,-1318,3218,-1234 $DEVICE_ID=1001
MM21 16 13 50 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=1916  $PIN_XY=3110,1832,3080,1916,3050,1832 $DEVICE_ID=1001
MM22 18 13 49 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=1454  $PIN_XY=3110,1538,3080,1454,3050,1538 $DEVICE_ID=1001
MM23 14 13 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=992  $PIN_XY=3110,908,3080,992,3050,908 $DEVICE_ID=1001
MM24 27 13 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=530  $PIN_XY=3110,614,3080,530,3050,614 $DEVICE_ID=1001
MM25 17 13 48 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=68  $PIN_XY=3110,-16,3080,68,3050,-16 $DEVICE_ID=1001
MM26 15 13 47 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=-394  $PIN_XY=3110,-310,3080,-394,3050,-310 $DEVICE_ID=1001
MM27 29 13 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=-856  $PIN_XY=3110,-940,3080,-856,3050,-940 $DEVICE_ID=1001
MM28 28 13 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=-1318  $PIN_XY=3110,-1234,3080,-1318,3050,-1234 $DEVICE_ID=1001
MM29 50 11 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=1916  $PIN_XY=2942,1832,2912,1916,2882,1832 $DEVICE_ID=1001
MM30 49 7 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=1475  $PIN_XY=2942,1538,2912,1475,2882,1538 $DEVICE_ID=1001
MM31 48 9 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=47  $PIN_XY=2942,-16,2912,47,2882,-16 $DEVICE_ID=1001
MM32 47 6 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=-373  $PIN_XY=2942,-310,2912,-373,2882,-310 $DEVICE_ID=1001
MM33 13 WEN GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2408 $Y=992  $PIN_XY=2438,908,2408,992,2378,908 $DEVICE_ID=1001
MM34 GND! 5 10 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2072 $Y=1454  $PIN_XY=2102,1538,2072,1454,2042,1538 $DEVICE_ID=1001
MM35 GND! 4 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2072 $Y=-394  $PIN_XY=2102,-310,2072,-394,2042,-310 $DEVICE_ID=1001
MM36 11 7 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1904 $Y=1937  $PIN_XY=1934,1832,1904,1937,1874,1832 $DEVICE_ID=1001
MM37 9 6 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1904 $Y=68  $PIN_XY=1934,-16,1904,68,1874,-16 $DEVICE_ID=1001
MM38 7 32 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1400 $Y=1916  $PIN_XY=1430,1832,1400,1916,1370,1832 $DEVICE_ID=1001
MM39 6 45 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1400 $Y=47  $PIN_XY=1430,-16,1400,47,1370,-16 $DEVICE_ID=1001
MM40 32 33 46 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=896 $Y=1916  $PIN_XY=926,1832,896,1916,866,1832 $DEVICE_ID=1001
MM41 45 43 44 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=896 $Y=47  $PIN_XY=926,-16,896,47,866,-16 $DEVICE_ID=1001
MM42 46 A0 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=728 $Y=1916  $PIN_XY=758,1832,728,1916,698,1832 $DEVICE_ID=1001
MM43 44 A1 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=728 $Y=47  $PIN_XY=758,-16,728,47,698,-16 $DEVICE_ID=1001
MM44 33 WEN GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=224 $Y=1937  $PIN_XY=254,1832,224,1937,194,1832 $DEVICE_ID=1001
MM45 43 WEN GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=224 $Y=68  $PIN_XY=254,-16,224,68,194,-16 $DEVICE_ID=1001
MM46 VDD! 16 WS0BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=2017  $PIN_XY=4118,2002,4088,2017,4058,2002 $DEVICE_ID=1003
MM47 VDD! 18 WS0 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=1353  $PIN_XY=4118,1368,4088,1353,4058,1368 $DEVICE_ID=1003
MM48 VDD! 14 RS0BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=1093  $PIN_XY=4118,1078,4088,1093,4058,1078 $DEVICE_ID=1003
MM49 VDD! 27 RS0 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=429  $PIN_XY=4118,444,4088,429,4058,444 $DEVICE_ID=1003
MM50 VDD! 17 WS1BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=169  $PIN_XY=4118,154,4088,169,4058,154 $DEVICE_ID=1003
MM51 VDD! 15 WS1 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=-495  $PIN_XY=4118,-480,4088,-495,4058,-480 $DEVICE_ID=1003
MM52 VDD! 29 RS1BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=-755  $PIN_XY=4118,-770,4088,-755,4058,-770 $DEVICE_ID=1003
MM53 VDD! 28 RS1 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4088 $Y=-1419  $PIN_XY=4118,-1404,4088,-1419,4058,-1404 $DEVICE_ID=1003
MM54 WS0BAR 16 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=2017  $PIN_XY=3950,2002,3920,2017,3890,2002 $DEVICE_ID=1003
MM55 WS0 18 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=1353  $PIN_XY=3950,1368,3920,1353,3890,1368 $DEVICE_ID=1003
MM56 RS0BAR 14 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=1093  $PIN_XY=3950,1078,3920,1093,3890,1078 $DEVICE_ID=1003
MM57 RS0 27 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=429  $PIN_XY=3950,444,3920,429,3890,444 $DEVICE_ID=1003
MM58 WS1BAR 17 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=169  $PIN_XY=3950,154,3920,169,3890,154 $DEVICE_ID=1003
MM59 WS1 15 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=-495  $PIN_XY=3950,-480,3920,-495,3890,-480 $DEVICE_ID=1003
MM60 RS1BAR 29 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=-755  $PIN_XY=3950,-770,3920,-755,3890,-770 $DEVICE_ID=1003
MM61 RS1 28 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3920 $Y=-1419  $PIN_XY=3950,-1404,3920,-1419,3890,-1404 $DEVICE_ID=1003
MM62 VDD! 16 WS0BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=1916  $PIN_XY=3782,2002,3752,1916,3722,2002 $DEVICE_ID=1003
MM63 VDD! 18 WS0 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=1454  $PIN_XY=3782,1368,3752,1454,3722,1368 $DEVICE_ID=1003
MM64 VDD! 14 RS0BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=992  $PIN_XY=3782,1078,3752,992,3722,1078 $DEVICE_ID=1003
MM65 VDD! 27 RS0 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=530  $PIN_XY=3782,444,3752,530,3722,444 $DEVICE_ID=1003
MM66 VDD! 17 WS1BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=68  $PIN_XY=3782,154,3752,68,3722,154 $DEVICE_ID=1003
MM67 VDD! 15 WS1 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=-394  $PIN_XY=3782,-480,3752,-394,3722,-480 $DEVICE_ID=1003
MM68 VDD! 29 RS1BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=-856  $PIN_XY=3782,-770,3752,-856,3722,-770 $DEVICE_ID=1003
MM69 VDD! 28 RS1 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3752 $Y=-1318  $PIN_XY=3782,-1404,3752,-1318,3722,-1404 $DEVICE_ID=1003
MM70 WS0BAR 16 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=1916  $PIN_XY=3614,2002,3584,1916,3554,2002 $DEVICE_ID=1003
MM71 WS0 18 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=1454  $PIN_XY=3614,1368,3584,1454,3554,1368 $DEVICE_ID=1003
MM72 RS0BAR 14 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=992  $PIN_XY=3614,1078,3584,992,3554,1078 $DEVICE_ID=1003
MM73 RS0 27 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=530  $PIN_XY=3614,444,3584,530,3554,444 $DEVICE_ID=1003
MM74 WS1BAR 17 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=68  $PIN_XY=3614,154,3584,68,3554,154 $DEVICE_ID=1003
MM75 WS1 15 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-394  $PIN_XY=3614,-480,3584,-394,3554,-480 $DEVICE_ID=1003
MM76 RS1BAR 29 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-856  $PIN_XY=3614,-770,3584,-856,3554,-770 $DEVICE_ID=1003
MM77 RS1 28 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3584 $Y=-1318  $PIN_XY=3614,-1404,3584,-1318,3554,-1404 $DEVICE_ID=1003
MM78 VDD! 5 56 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=971  $PIN_XY=3278,1078,3248,971,3218,1078 $DEVICE_ID=1003
MM79 VDD! 10 55 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=551  $PIN_XY=3278,444,3248,551,3218,444 $DEVICE_ID=1003
MM80 VDD! 4 53 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=-877  $PIN_XY=3278,-770,3248,-877,3218,-770 $DEVICE_ID=1003
MM81 VDD! 8 54 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3248 $Y=-1318  $PIN_XY=3278,-1404,3248,-1318,3218,-1404 $DEVICE_ID=1003
MM82 VDD! 13 16 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=1916  $PIN_XY=3110,2002,3080,1916,3050,2002 $DEVICE_ID=1003
MM83 VDD! 13 18 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=1454  $PIN_XY=3110,1368,3080,1454,3050,1368 $DEVICE_ID=1003
MM84 56 13 14 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=992  $PIN_XY=3110,1078,3080,992,3050,1078 $DEVICE_ID=1003
MM85 55 13 27 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=530  $PIN_XY=3110,444,3080,530,3050,444 $DEVICE_ID=1003
MM86 VDD! 13 17 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=68  $PIN_XY=3110,154,3080,68,3050,154 $DEVICE_ID=1003
MM87 VDD! 13 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3080 $Y=-394  $PIN_XY=3110,-480,3080,-394,3050,-480 $DEVICE_ID=1003
MM88 53 13 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=-856  $PIN_XY=3110,-770,3080,-856,3050,-770 $DEVICE_ID=1003
MM89 54 13 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3080 $Y=-1318  $PIN_XY=3110,-1404,3080,-1318,3050,-1404 $DEVICE_ID=1003
MM90 16 11 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=1916  $PIN_XY=2942,2002,2912,1916,2882,2002 $DEVICE_ID=1003
MM91 18 7 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=1475  $PIN_XY=2942,1368,2912,1475,2882,1368 $DEVICE_ID=1003
MM92 17 9 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=47  $PIN_XY=2942,154,2912,47,2882,154 $DEVICE_ID=1003
MM93 15 6 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2912 $Y=-373  $PIN_XY=2942,-480,2912,-373,2882,-480 $DEVICE_ID=1003
MM94 VDD! WEN 13 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2576 $Y=1072  $PIN_XY=2606,1078,2576,1072,2546,1078 $DEVICE_ID=1003
MM95 13 WEN VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2408 $Y=992  $PIN_XY=2438,1078,2408,992,2378,1078 $DEVICE_ID=1003
MM96 VDD! 7 11 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2072 $Y=2017  $PIN_XY=2102,2002,2072,2017,2042,2002 $DEVICE_ID=1003
MM97 VDD! 5 10 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2072 $Y=1454  $PIN_XY=2102,1368,2072,1454,2042,1368 $DEVICE_ID=1003
MM98 VDD! 6 9 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2072 $Y=154  $PIN_XY=2102,154,2072,154,2042,154 $DEVICE_ID=1003
MM99 VDD! 4 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2072 $Y=-394  $PIN_XY=2102,-480,2072,-394,2042,-480 $DEVICE_ID=1003
MM100 11 7 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1904 $Y=1937  $PIN_XY=1934,2002,1904,1937,1874,2002 $DEVICE_ID=1003
MM101 10 5 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1904 $Y=1374  $PIN_XY=1934,1368,1904,1374,1874,1368 $DEVICE_ID=1003
MM102 9 6 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1904 $Y=68  $PIN_XY=1934,154,1904,68,1874,154 $DEVICE_ID=1003
MM103 8 4 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1904 $Y=-474  $PIN_XY=1934,-480,1904,-474,1874,-480 $DEVICE_ID=1003
MM104 VDD! 32 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1568 $Y=2017  $PIN_XY=1598,2002,1568,2017,1538,2002 $DEVICE_ID=1003
MM105 VDD! 52 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1568 $Y=1374  $PIN_XY=1598,1368,1568,1374,1538,1368 $DEVICE_ID=1003
MM106 VDD! 45 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1568 $Y=148  $PIN_XY=1598,154,1568,148,1538,154 $DEVICE_ID=1003
MM107 VDD! 51 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1568 $Y=-474  $PIN_XY=1598,-480,1568,-474,1538,-480 $DEVICE_ID=1003
MM108 7 32 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1400 $Y=1916  $PIN_XY=1430,2002,1400,1916,1370,2002 $DEVICE_ID=1003
MM109 5 52 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1400 $Y=1475  $PIN_XY=1430,1368,1400,1475,1370,1368 $DEVICE_ID=1003
MM110 6 45 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1400 $Y=47  $PIN_XY=1430,154,1400,47,1370,154 $DEVICE_ID=1003
MM111 4 51 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1400 $Y=-373  $PIN_XY=1430,-480,1400,-373,1370,-480 $DEVICE_ID=1003
MM112 VDD! 33 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=896 $Y=1916  $PIN_XY=926,2002,896,1916,866,2002 $DEVICE_ID=1003
MM113 VDD! WEN 52 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=896 $Y=1475  $PIN_XY=926,1368,896,1475,866,1368 $DEVICE_ID=1003
MM114 VDD! 43 45 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=896 $Y=47  $PIN_XY=926,154,896,47,866,154 $DEVICE_ID=1003
MM115 VDD! WEN 51 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=896 $Y=-373  $PIN_XY=926,-480,896,-373,866,-480 $DEVICE_ID=1003
MM116 32 A0 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=728 $Y=1916  $PIN_XY=758,2002,728,1916,698,2002 $DEVICE_ID=1003
MM117 52 A0 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=728 $Y=1475  $PIN_XY=758,1368,728,1475,698,1368 $DEVICE_ID=1003
MM118 45 A1 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=728 $Y=47  $PIN_XY=758,154,728,47,698,154 $DEVICE_ID=1003
MM119 51 A1 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=728 $Y=-373  $PIN_XY=758,-480,728,-373,698,-480 $DEVICE_ID=1003
MM120 VDD! WEN 33 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=392 $Y=2017  $PIN_XY=422,2002,392,2017,362,2002 $DEVICE_ID=1003
MM121 VDD! WEN 43 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=392 $Y=148  $PIN_XY=422,154,392,148,362,154 $DEVICE_ID=1003
MM122 33 WEN VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=224 $Y=1937  $PIN_XY=254,2002,224,1937,194,2002 $DEVICE_ID=1003
MM123 43 WEN VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=224 $Y=68  $PIN_XY=254,154,224,68,194,154 $DEVICE_ID=1003
XXCE9F2C661 GND! VDD! 8 4 36 39 inv $T=2294 -100 0 180 $X=1682 $Y=-690
XXCE9F2C662 GND! VDD! 9 6 36 40 inv $T=1682 -226 0 0 $X=1682 $Y=-226
XXCE9F2C663 GND! VDD! 13 WEN 35 41 inv $T=2186 698 0 0 $X=2186 $Y=698
XXCE9F2C664 GND! VDD! 10 5 37 41 inv $T=2294 1748 0 180 $X=1682 $Y=1158
XXCE9F2C665 GND! VDD! 11 7 37 42 inv $T=1682 1622 0 0 $X=1682 $Y=1622
XXCE9F2C666 GND! VDD! _GENERATED_78 _GENERATED_77 34 38 sram_filler $T=4650 -1024 0 180 $X=4202 $Y=-1613
XXCE9F2C667 GND! VDD! _GENERATED_80 _GENERATED_79 34 39 sram_filler $T=4198 -1150 0 0 $X=4202 $Y=-1150
XXCE9F2C668 GND! VDD! _GENERATED_82 _GENERATED_81 36 39 sram_filler $T=4650 -100 0 180 $X=4202 $Y=-690
XXCE9F2C669 GND! VDD! _GENERATED_84 _GENERATED_83 36 40 sram_filler $T=4198 -226 0 0 $X=4202 $Y=-226
XXCE9F2C6610 GND! VDD! _GENERATED_86 _GENERATED_85 35 40 sram_filler $T=4650 824 0 180 $X=4202 $Y=234
XXCE9F2C6611 GND! VDD! _GENERATED_88 _GENERATED_87 35 41 sram_filler $T=4198 698 0 0 $X=4202 $Y=698
XXCE9F2C6612 GND! VDD! _GENERATED_90 _GENERATED_89 37 41 sram_filler $T=4650 1748 0 180 $X=4202 $Y=1158
XXCE9F2C6613 GND! VDD! _GENERATED_92 _GENERATED_91 37 42 sram_filler $T=4198 1622 0 0 $X=4202 $Y=1622
XXCE9F2C6614 GND! VDD! _GENERATED_94 _GENERATED_93 34 38 sram_filler $T=-2 -1024 1 0 $X=2 $Y=-1613
XXCE9F2C6615 GND! VDD! _GENERATED_95 GND! 34 38 sram_filler $T=334 -1024 1 0 $X=338 $Y=-1613
XXCE9F2C6616 GND! VDD! VDD! _GENERATED_96 34 38 sram_filler $T=502 -1024 1 0 $X=506 $Y=-1613
XXCE9F2C6617 GND! VDD! _GENERATED_97 GND! 34 39 sram_filler $T=-2 -1150 0 0 $X=2 $Y=-1150
XXCE9F2C6618 GND! VDD! VDD! _GENERATED_98 34 39 sram_filler $T=166 -1150 0 0 $X=170 $Y=-1150
XXCE9F2C6619 GND! VDD! _GENERATED_100 _GENERATED_99 34 39 sram_filler $T=502 -1150 0 0 $X=506 $Y=-1150
XXCE9F2C6620 GND! VDD! VDD! _GENERATED_101 34 38 sram_filler $T=1342 -1024 1 0 $X=1346 $Y=-1613
XXCE9F2C6621 GND! VDD! _GENERATED_102 GND! 34 38 sram_filler $T=1174 -1024 1 0 $X=1178 $Y=-1613
XXCE9F2C6622 GND! VDD! _GENERATED_104 _GENERATED_103 34 38 sram_filler $T=838 -1024 1 0 $X=842 $Y=-1613
XXCE9F2C6623 GND! VDD! VDD! _GENERATED_105 34 39 sram_filler $T=1342 -1150 0 0 $X=1346 $Y=-1150
XXCE9F2C6624 GND! VDD! _GENERATED_106 GND! 34 39 sram_filler $T=1174 -1150 0 0 $X=1178 $Y=-1150
XXCE9F2C6625 GND! VDD! _GENERATED_108 _GENERATED_107 34 39 sram_filler $T=838 -1150 0 0 $X=842 $Y=-1150
XXCE9F2C6626 GND! VDD! _GENERATED_110 _GENERATED_109 34 39 sram_filler $T=1678 -1150 0 0 $X=1682 $Y=-1150
XXCE9F2C6627 GND! VDD! _GENERATED_112 _GENERATED_111 34 38 sram_filler $T=2130 -1024 0 180 $X=1682 $Y=-1613
XXCE9F2C6628 GND! VDD! VDD! _GENERATED_113 35 41 sram_filler $T=1846 698 0 0 $X=1850 $Y=698
XXCE9F2C6629 GND! VDD! _GENERATED_114 GND! 35 40 sram_filler $T=2298 824 0 180 $X=1850 $Y=234
XXCE9F2C6630 GND! VDD! _GENERATED_116 _GENERATED_115 34 39 sram_filler $T=2014 -1150 0 0 $X=2018 $Y=-1150
XXCE9F2C6631 GND! VDD! _GENERATED_118 _GENERATED_117 34 38 sram_filler $T=2466 -1024 0 180 $X=2018 $Y=-1613
XXCE9F2C6632 GND! VDD! _GENERATED_120 _GENERATED_119 34 38 sram_filler $T=2802 -1024 0 180 $X=2354 $Y=-1613
XXCE9F2C6633 GND! VDD! _GENERATED_122 _GENERATED_121 34 39 sram_filler $T=2350 -1150 0 0 $X=2354 $Y=-1150
XXCE9F2C6634 GND! VDD! _GENERATED_124 _GENERATED_123 35 40 sram_filler $T=1794 824 0 180 $X=1346 $Y=234
XXCE9F2C6635 GND! VDD! _GENERATED_126 _GENERATED_125 35 40 sram_filler $T=1458 824 0 180 $X=1010 $Y=234
XXCE9F2C6636 GND! VDD! _GENERATED_128 _GENERATED_127 35 40 sram_filler $T=1122 824 0 180 $X=674 $Y=234
XXCE9F2C6637 GND! VDD! _GENERATED_130 _GENERATED_129 35 40 sram_filler $T=786 824 0 180 $X=338 $Y=234
XXCE9F2C6638 GND! VDD! _GENERATED_132 _GENERATED_131 35 40 sram_filler $T=450 824 0 180 $X=2 $Y=234
XXCE9F2C6639 GND! VDD! VDD! _GENERATED_133 35 41 sram_filler $T=1342 698 0 0 $X=1346 $Y=698
XXCE9F2C6640 GND! VDD! _GENERATED_134 GND! 35 41 sram_filler $T=1174 698 0 0 $X=1178 $Y=698
XXCE9F2C6641 GND! VDD! _GENERATED_136 _GENERATED_135 35 41 sram_filler $T=838 698 0 0 $X=842 $Y=698
XXCE9F2C6642 GND! VDD! VDD! _GENERATED_137 35 41 sram_filler $T=502 698 0 0 $X=506 $Y=698
XXCE9F2C6643 GND! VDD! _GENERATED_138 GND! 35 41 sram_filler $T=334 698 0 0 $X=338 $Y=698
XXCE9F2C6644 GND! VDD! _GENERATED_140 _GENERATED_139 35 41 sram_filler $T=-2 698 0 0 $X=2 $Y=698
XXCE9F2C6645 GND! VDD! _GENERATED_141 GND! 36 39 sram_filler $T=2802 -100 0 180 $X=2354 $Y=-690
XXCE9F2C6646 GND! VDD! VDD! _GENERATED_142 36 39 sram_filler $T=2634 -100 0 180 $X=2186 $Y=-690
XXCE9F2C6647 GND! VDD! _GENERATED_143 GND! 36 40 sram_filler $T=2182 -226 0 0 $X=2186 $Y=-226
XXCE9F2C6648 GND! VDD! VDD! _GENERATED_144 36 40 sram_filler $T=2350 -226 0 0 $X=2354 $Y=-226
XXCE9F2C6649 GND! VDD! _GENERATED_145 GND! 35 40 sram_filler $T=2802 824 0 180 $X=2354 $Y=234
XXCE9F2C6650 GND! VDD! VDD! _GENERATED_146 35 40 sram_filler $T=2634 824 0 180 $X=2186 $Y=234
XXCE9F2C6651 GND! VDD! _GENERATED_147 GND! 37 41 sram_filler $T=2802 1748 0 180 $X=2354 $Y=1158
XXCE9F2C6652 GND! VDD! VDD! _GENERATED_148 37 41 sram_filler $T=2634 1748 0 180 $X=2186 $Y=1158
XXCE9F2C6653 GND! VDD! VDD! _GENERATED_149 37 42 sram_filler $T=2350 1622 0 0 $X=2354 $Y=1622
XXCE9F2C6654 GND! VDD! _GENERATED_150 GND! 37 42 sram_filler $T=2182 1622 0 0 $X=2186 $Y=1622
XXCE9F2C6655 GND! VDD! _GENERATED_151 GND! 35 41 sram_filler $T=1678 698 0 0 $X=1682 $Y=698
XXCE9F2C6656 GND! VDD! VDD! _GENERATED_152 35 40 sram_filler $T=2130 824 0 180 $X=1682 $Y=234
XXCE9F2C6657 GND! VDD! WS1BAR 17 15 27 15 27 27 27 36 
+	40 invx4 $T=3338 -226 0 0 $X=3362 $Y=-226
XXCE9F2C6658 GND! VDD! RS0 27 14 17 14 17 17 17 35 
+	40 invx4 $T=3338 824 1 0 $X=3362 $Y=234
XXCE9F2C6659 GND! VDD! RS1 28 29 69 29 71 73 75 34 
+	38 invx4 $T=3338 -1024 1 0 $X=3362 $Y=-1613
XXCE9F2C6660 GND! VDD! WS1 15 17 29 17 29 29 29 36 
+	39 invx4 $T=3338 -100 1 0 $X=3362 $Y=-690
XXCE9F2C6661 GND! VDD! RS1BAR 29 28 15 28 15 15 15 34 
+	39 invx4 $T=3338 -1150 0 0 $X=3362 $Y=-1150
XXCE9F2C6662 GND! VDD! WS0BAR 16 18 70 18 72 74 76 37 
+	42 invx4 $T=3338 1622 0 0 $X=3362 $Y=1622
XXCE9F2C6663 GND! VDD! WS0 18 16 14 16 14 14 14 37 
+	41 invx4 $T=3338 1748 1 0 $X=3362 $Y=1158
XXCE9F2C6664 GND! VDD! RS0BAR 14 27 18 27 18 18 18 35 
+	41 invx4 $T=3338 698 0 0 $X=3362 $Y=698
XXCE9F2C6665 GND! VDD! VDD! WEN 43 A1 51 45 4 6 36 
+	40 39 44 Demux $T=2 -688 0 0 $X=2 $Y=-690
XXCE9F2C6666 GND! VDD! VDD! WEN 33 A0 52 32 5 7 37 
+	42 41 46 Demux $T=2 1160 0 0 $X=2 $Y=1158
XXCE9F2C6667 GND! VDD! 15 6 13 9 13 47 36 39 nand $T=2272 128 1 0 $X=2690 $Y=-690
XXCE9F2C6668 GND! VDD! 17 9 13 6 13 48 36 40 nand $T=2272 -454 0 0 $X=2690 $Y=-226
XXCE9F2C6669 GND! VDD! 18 7 13 11 13 49 37 41 nand $T=2272 1976 1 0 $X=2690 $Y=1158
XXCE9F2C6670 GND! VDD! 16 11 13 7 13 50 37 42 nand $T=2272 1394 0 0 $X=2690 $Y=1622
XXCE9F2C6671 GND! VDD! 29 4 13 8 13 13 53 34 39 nor $T=4098 -1152 1 180 $X=2690 $Y=-1150
XXCE9F2C6672 GND! VDD! 28 8 13 4 13 68 54 34 38 nor $T=4098 -1022 0 180 $X=2690 $Y=-1613
XXCE9F2C6673 GND! VDD! 27 10 13 5 13 13 55 35 40 nor $T=4098 826 0 180 $X=2690 $Y=234
XXCE9F2C6674 GND! VDD! 14 5 13 10 13 13 56 35 41 nor $T=4098 696 1 180 $X=2690 $Y=698
.ends agen_unit
