*  Generated for: PrimeSim
*  Design library name: group8
*  Design cell name: tb2025_2_tree_decoder
*  Design view name: schematic
.option search='/mnt/designkits/ncsu/FreePDK3/hspice/models'

.param clkperiod=90p clkrise=5p vdd=0.8
.option PARHIER = LOCAL
.include '/mnt/coe/workspace/ece/ece546-spr25/group8/group8_project/invec.dat'

.include '/mnt/coe/workspace/ece/ece546-spr25/group8/group8_project/outvec.dat'
.option PORT_VOLTAGE_SCALE_TO_2X = 1
.option S_ELEM_CACHE_DIR = "/mnt/ncsudrive/n/nbandeh/.synopsys_custom/sparam_dir"
.option PVA_OUTPUT_DIR = "/mnt/ncsudrive/n/nbandeh/.synopsys_custom/pva_dir"

.option WDF=1
.temp 25
.lib 'fet.mod' nfet_typ
.lib 'fet.mod' pfet_typ

*PrimeWave Design Environment Based on Custom Infrastructure
*Version W-2024.09-SP1-2
*Thu Apr 10 17:21:14 2025

.global gnd! vdd!
********************************************************************************
* Library          : proj_common
* Cell             : inputbuf
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt inputbuf out in
m9 out net7 gnd! nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m8 net7 in gnd! nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m12 net7 in vdd! pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m13 out net7 vdd! pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
.ends inputbuf

********************************************************************************
* Library          : group8
* Cell             : precharge_logic
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt precharge_logic bl bl_bar clk
m5 bl_bar clk vdd! pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m4 vdd! clk bl pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m3 bl clk bl_bar pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
.ends precharge_logic

********************************************************************************
* Library          : group8
* Cell             : sram_6t
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt sram_6t bl bl_bar wl
m1 qbar q vdd! pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
m0 q qbar vdd! pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
m5 bl wl q nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
m6 qbar wl bl_bar nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
m3 qbar q gnd! nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
m2 q qbar gnd! nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
.ends sram_6t

********************************************************************************
* Library          : group8
* Cell             : nand
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt nand a b y
m1 net4 b gnd! nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m0 y a net4 nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m3 y b vdd! pfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
m2 y a vdd! pfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
.ends nand

********************************************************************************
* Library          : group8
* Cell             : inv
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt inv in out
m0 out in vdd! pfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
m1 out in gnd! nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=1.17e-07 pseo=1.17e-07
.ends inv

********************************************************************************
* Library          : group8
* Cell             : buffer_highdrive
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt buffer_highdrive in out
m4 net9 in vdd! pfet nfin=8 adeo=2.268e-15 aseo=2.268e-15 pdeo=4.68e-07 pseo=4.68e-07
m0 out net9 vdd! pfet nfin=20 adeo=5.67e-15 aseo=5.67e-15 pdeo=1.17e-06 pseo=1.17e-06
m5 net9 in gnd! nfet nfin=8 adeo=2.268e-15 aseo=2.268e-15 pdeo=4.68e-07 pseo=4.68e-07
m1 out net9 gnd! nfet nfin=20 adeo=5.67e-15 aseo=5.67e-15 pdeo=1.17e-06 pseo=1.17e-06
.ends buffer_highdrive

********************************************************************************
* Library          : group8
* Cell             : invx4
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt invx4 in out
m0 out in vdd! pfet nfin=8 adeo=2.268e-15 aseo=2.268e-15 pdeo=4.68e-07 pseo=4.68e-07
m1 out in gnd! nfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
.ends invx4

********************************************************************************
* Library          : group8
* Cell             : nor
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt nor a b y
m1 y b gnd! nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m0 y a gnd! nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m3 net11 a vdd! pfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
m2 y b net11 pfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
.ends nor

********************************************************************************
* Library          : group8
* Cell             : static_row_decoder_3by8
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt static_row_decoder_3by8 a0 a1 a2 wlref y0 y1 y2 y3 y4 y5 y6 y7
xi107 a2 a1 net176 nand
xi106 a0 net181 net177 nand
xi104 a2 a1 net169 nand
xi103 net173 net181 net170 nand
xi101 a2 net182 net162 nand
xi100 a0 net181 net163 nand
xi98 a2 net182 net155 nand
xi97 net173 net181 net156 nand
xi95 net121 a1 net148 nand
xi94 a0 net181 net149 nand
xi86 net121 net181 net132 nand
xi85 net173 net182 net131 nand
xi89 net121 net182 net134 nand
xi91 net173 net181 net142 nand
xi92 net121 a1 net141 nand
xi88 a0 net181 net135 nand
xi83 a2 net121 inv
xi82 net130 y0 buffer_highdrive
xi80 net133 y1 buffer_highdrive
xi79 net140 y2 buffer_highdrive
xi78 net147 y3 buffer_highdrive
xi77 net154 y4 buffer_highdrive
xi76 net161 y5 buffer_highdrive
xi75 net168 y6 buffer_highdrive
xi74 net175 y7 buffer_highdrive
xi109 wlref net181 buffer_highdrive
xi18 a0 net173 invx4
xi17 a1 net182 invx4
xi108 net176 net177 net175 nor
xi105 net169 net170 net168 nor
xi102 net162 net163 net161 nor
xi99 net155 net156 net154 nor
xi96 net148 net149 net147 nor
xi87 net131 net132 net130 nor
xi90 net134 net135 net133 nor
xi93 net141 net142 net140 nor
.ends static_row_decoder_3by8

********************************************************************************
* Library          : group8
* Cell             : 2to4_decoder
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt _2to4_decoder bl0 bl0_bar bl1 bl1_bar bl2 bl2_bar bl3 bl3_bar in0 in0bar
+  op0 op0bar rs0 rs0bar rs1 rs1bar ws0 ws0bar ws1 ws1bar
m53 op0 rs1 rd23 pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m52 op0bar rs1 rdb23 pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m51 op0 rs1bar rd01 pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m50 op0bar rs1bar rdb01 pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m49 rdb01 rs0bar bl0_bar pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m48 rd23 rs0 bl3 pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m47 rdb23 rs0 bl3_bar pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m46 rd23 rs0bar bl2 pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m45 rdb23 rs0bar bl2_bar pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m44 rd01 rs0 bl1 pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m43 rdb01 rs0 bl1_bar pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m42 rd01 rs0bar bl0 pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m31 bl0 ws0bar wd01 nfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07
+ pseo=2.34e-07
m30 bl0_bar ws0bar wdb01 nfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07
+  pseo=2.34e-07
m41 wd23 ws1 in0 nfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
m40 wdb23 ws1 in0bar nfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07
+ pseo=2.34e-07
m39 wd01 ws1bar in0 nfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07
+ pseo=2.34e-07
m38 wdb01 ws1bar in0bar nfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07
+ pseo=2.34e-07
m37 bl3 ws0 wd23 nfet nfin=6 adeo=1.701e-15 aseo=1.701e-15 pdeo=3.51e-07 pseo=3.51e-07
m36 bl3_bar ws0 wdb23 nfet nfin=6 adeo=1.701e-15 aseo=1.701e-15 pdeo=3.51e-07
+ pseo=3.51e-07
m35 bl2 ws0bar wd23 nfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07
+ pseo=2.34e-07
m34 bl2_bar ws0bar wdb23 nfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07
+  pseo=2.34e-07
m33 bl1 ws0 wd01 nfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
m32 bl1_bar ws0 wdb01 nfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07
+ pseo=2.34e-07
.ends _2to4_decoder

********************************************************************************
* Library          : group8
* Cell             : columnDecoder
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt columndecoder bl0 bl0bar bl1 bl1bar bl2 bl2bar bl3 bl3bar bl4 bl4bar bl5
+  bl5bar bl6 bl6bar bl7 bl7bar bl8 bl8bar bl9 bl9bar bl10 bl10bar bl11 bl11bar
+ bl12 bl12bar bl13 bl13bar bl14 bl14bar bl15 bl15bar i0 i0bar i1 i1bar i2 i2bar
+  i3 i3bar q0 q0baar q1 q1bar q2 q2bar q3 q3bar rs0 rs0bar rs1 rs1bar ws0
+ ws0bar ws1 ws1bar
xi3 bl12 bl12bar bl13 bl13bar bl14 bl14bar bl15 bl15bar i3 i3bar q3 q3bar rs0
+ rs0bar rs1 rs1bar ws0 ws0bar ws1 ws1bar _2to4_decoder
xi2 bl8 bl8bar bl9 bl9bar bl10 bl10bar bl11 bl11bar i2 i2bar q2 q2bar rs0 rs0bar
+ rs1 rs1bar ws0 ws0bar ws1 ws1bar _2to4_decoder
xi1 bl4 bl4bar bl5 bl5bar bl6 bl6bar bl7 bl7bar i1 i1bar q1 q1bar rs0 rs0bar rs1
+ rs1bar ws0 ws0bar ws1 ws1bar _2to4_decoder
xi0 bl0 bl0bar bl1 bl1bar bl2 bl2bar bl3bar bl3 i0 i0bar q0 q0baar rs0 rs0bar
+ rs1 rs1bar ws0 ws0bar ws1 ws1bar _2to4_decoder
.ends columndecoder

********************************************************************************
* Library          : group8
* Cell             : Write_Driver
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt write_driver din wbdata wdata
m18 net33 din vdd! pfet nfin=8 adeo=2.268e-15 aseo=2.268e-15 pdeo=4.68e-07 pseo=4.68e-07
m13 net26 din vdd! pfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
m12 net25 net26 vdd! pfet nfin=8 adeo=2.268e-15 aseo=2.268e-15 pdeo=4.68e-07
+ pseo=4.68e-07
m17 net32 net33 vdd! pfet nfin=16 adeo=4.536e-15 aseo=4.536e-15 pdeo=9.36e-07
+ pseo=9.36e-07
m16 wbdata net32 vdd! pfet nfin=20 adeo=5.67e-15 aseo=5.67e-15 pdeo=1.17e-06
+ pseo=1.17e-06
m1 wdata net35 vdd! pfet nfin=20 adeo=5.67e-15 aseo=5.67e-15 pdeo=1.17e-06 pseo=1.17e-06
m0 net35 net25 vdd! pfet nfin=16 adeo=4.536e-15 aseo=4.536e-15 pdeo=9.36e-07
+ pseo=9.36e-07
m21 net33 din gnd! nfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07 pseo=2.34e-07
m20 net32 net33 gnd! nfet nfin=8 adeo=2.268e-15 aseo=2.268e-15 pdeo=4.68e-07
+ pseo=4.68e-07
m19 wbdata net32 gnd! nfet nfin=10 adeo=2.835e-15 aseo=2.835e-15 pdeo=5.85e-07
+ pseo=5.85e-07
m15 net26 din gnd! nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m14 net25 net26 gnd! nfet nfin=4 adeo=1.134e-15 aseo=1.134e-15 pdeo=2.34e-07
+ pseo=2.34e-07
m5 wdata net35 gnd! nfet nfin=10 adeo=2.835e-15 aseo=2.835e-15 pdeo=5.85e-07
+ pseo=5.85e-07
m4 net35 net25 gnd! nfet nfin=8 adeo=2.268e-15 aseo=2.268e-15 pdeo=4.68e-07
+ pseo=4.68e-07
.ends write_driver

********************************************************************************
* Library          : group8
* Cell             : read_circuit
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt read_circuit bl blbar out
xi0 bl net6 net2 nand
xi1 net2 out inv
xi2 blbar net6 invx4
.ends read_circuit

********************************************************************************
* Library          : group8
* Cell             : tspc_pos_ff
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt tspc_pos_ff d q phi
m16 q net26 gnd! nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m4 net26 phi net14 nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m3 net27 net17 net11 nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m2 net14 net27 gnd! nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m1 net11 phi gnd! nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m0 net17 d gnd! nfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m15 q net26 vdd! pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m8 net26 net27 vdd! pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m7 net27 phi vdd! pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m6 net20 d vdd! pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
m5 net17 phi net20 pfet nfin=2 adeo=5.67e-16 aseo=5.67e-16 pdeo=117n pseo=117n
.ends tspc_pos_ff

********************************************************************************
* Library          : group8
* Cell             : Demux
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt demux a sel y0 y1
xi1 sel a net12 nand
xi0 net7 a net10 nand
xi4 net12 y1 inv
xi3 net10 y0 inv
xi2 sel net7 inv
.ends demux

********************************************************************************
* Library          : group8
* Cell             : agen_unit
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt agen_unit a0 a1 rs0 rs0bar rs1 rs1bar wen ws0 ws0bar ws1 ws1bar
xi1 a1 wen net82 net88 demux
xi0 a0 wen net77 net86 demux
xi34 wen net75 inv
xi17 net88 net87 inv
xi16 net82 net81 inv
xi14 net77 net79 inv
xi15 net86 net85 inv
xi18 net86 net75 net43 nor
xi19 net85 net75 net46 nor
xi20 net88 net75 net49 nor
xi21 net87 net75 net52 nor
xi25 net82 net75 net64 nand
xi24 net81 net75 net61 nand
xi22 net79 net75 net55 nand
xi23 net77 net75 net58 nand
xi33 net52 rs1 invx4
xi32 net49 rs1bar invx4
xi31 net64 ws1 invx4
xi30 net61 ws1bar invx4
xi29 net46 rs0 invx4
xi28 net43 rs0bar invx4
xi27 net58 ws0 invx4
xi26 net55 ws0bar invx4
.ends agen_unit

********************************************************************************
* Library          : group8
* Cell             : buffer
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt buffer in out
xi1 net4 out inv
xi0 in net4 inv
.ends buffer

********************************************************************************
* Library          : group8
* Cell             : WLRef_PC
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt wlref_pc clk pc rsnew wlref clk_dff
xi60 net126 clk_dff buffer
xi59 net127 net126 buffer
xi58 net128 net127 buffer
xi57 net129 net128 buffer
xi56 net124 net129 buffer
xi55 net123 net124 buffer
xi54 net122 net123 buffer
xi53 net121 net122 buffer
xi52 net118 net121 buffer
xi51 net116 net118 buffer
xi50 net115 net116 buffer
xi49 net114 net115 buffer
xi46 net108 net110 buffer
xi48 net111 net114 buffer
xi47 net110 net111 buffer
xi21 net108 net59 buffer
xi19 net39 net62 buffer
xi20 net61 net39 buffer
xi14 net62 net60 buffer
xi8 net60 net108 buffer
xi0 clk net61 buffer
xi29 net76 rsnew invx4
xi10 net21 pc invx4
xi16 net36 wlref invx4
xi42 net103 net100 inv
xi40 net104 net103 inv
xi39 net100 net97 inv
xi38 net101 net104 inv
xi37 net97 net95 inv
xi36 net96 net101 inv
xi35 net89 net96 inv
xi34 net72 net94 inv
xi33 net94 net89 inv
xi32 net85 net84 inv
xi31 net84 net83 inv
xi30 net83 net72 inv
xi27 net95 clk_inverted_delayed inv
xi26 net106 net85 inv
xi25 net68 net106 inv
xi23 clk clk_inverted inv
xi24 clk_inverted net68 inv
xi28 clk_inverted_delayed clk_inverted net76 nor
xi13 net59 net61 net21 nor
xi15 net61 net60 net36 nand
.ends wlref_pc

********************************************************************************
* Library          : group8
* Cell             : inv_highdrive
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt inv_highdrive in out
m4 out in vdd! pfet nfin=20 adeo=5.67e-15 aseo=5.67e-15 pdeo=1.17e-06 pseo=1.17e-06
m5 out in gnd! nfet nfin=20 adeo=5.67e-15 aseo=5.67e-15 pdeo=1.17e-06 pseo=1.17e-06
.ends inv_highdrive

********************************************************************************
* Library          : group8
* Cell             : memory_array
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt memory_array a<0> a<1> a<2> a<3> a<4> clk d<0> d<1> d<2> d<3> q<0> q<1>
+ q<2> q<3> wenb
xi182 net573 net557 pc precharge_logic
xi147 bl3bar bl3 pc precharge_logic
xi146 net579 net563 pc precharge_logic
xi145 net578 net562 pc precharge_logic
xi144 net577 net561 pc precharge_logic
xi143 bl2bar bl2 pc precharge_logic
xi142 net575 net559 pc precharge_logic
xi141 net588 net572 pc precharge_logic
xi140 net587 net571 pc precharge_logic
xi139 bl1bar bl1 pc precharge_logic
xi138 net585 net569 pc precharge_logic
xi137 net584 net568 pc precharge_logic
xi136 net583 net652 pc precharge_logic
xi135 bl0bar bl0 pc precharge_logic
xi134 net581 net565 pc precharge_logic
xi133 net574 net558 pc precharge_logic
xi199 net557 net573 net546 sram_6t
xi55 net569 net585 net546 sram_6t
xi54 net568 net584 net546 sram_6t
xi53 net652 net583 net546 sram_6t
xi52 bl0 bl0bar net546 sram_6t
xi47 bl1 bl1bar net550 sram_6t
xi51 net565 net581 net546 sram_6t
xi50 net558 net574 net546 sram_6t
xi64 net571 net587 net655 sram_6t
xi65 net572 net588 net655 sram_6t
xi66 net559 net575 net655 sram_6t
xi67 bl2 bl2bar net655 sram_6t
xi68 net561 net577 net655 sram_6t
xi69 net562 net578 net655 sram_6t
xi70 net563 net579 net655 sram_6t
xi71 bl3 bl3bar net655 sram_6t
xi72 net571 net587 net556 sram_6t
xi73 net571 net587 net555 sram_6t
xi74 net572 net588 net555 sram_6t
xi75 net559 net575 net555 sram_6t
xi76 bl2 bl2bar net555 sram_6t
xi77 net561 net577 net555 sram_6t
xi104 bl3 bl3bar net548 sram_6t
xi103 net563 net579 net548 sram_6t
xi102 net562 net578 net548 sram_6t
xi101 net561 net577 net548 sram_6t
xi100 bl2 bl2bar net548 sram_6t
xi99 net559 net575 net548 sram_6t
xi98 net572 net588 net548 sram_6t
xi97 net571 net587 net548 sram_6t
xi95 bl3 bl3bar net551 sram_6t
xi94 net563 net579 net551 sram_6t
xi93 net562 net578 net551 sram_6t
xi92 net561 net577 net551 sram_6t
xi91 bl2 bl2bar net551 sram_6t
xi90 net559 net575 net551 sram_6t
xi89 net572 net588 net551 sram_6t
xi88 net571 net587 net551 sram_6t
xi87 bl3 bl3bar net556 sram_6t
xi86 net563 net579 net556 sram_6t
xi85 net562 net578 net556 sram_6t
xi84 net561 net577 net556 sram_6t
xi83 bl2 bl2bar net556 sram_6t
xi82 net559 net575 net556 sram_6t
xi81 net572 net588 net556 sram_6t
xi80 bl3 bl3bar net555 sram_6t
xi79 net563 net579 net555 sram_6t
xi78 net562 net578 net555 sram_6t
xi117 net561 net577 net546 sram_6t
xi116 bl2 bl2bar net546 sram_6t
xi115 net559 net575 net546 sram_6t
xi114 net572 net588 net546 sram_6t
xi113 net571 net587 net546 sram_6t
xi112 net571 net587 net544 sram_6t
xi111 bl3 bl3bar net550 sram_6t
xi110 net563 net579 net550 sram_6t
xi109 net562 net578 net550 sram_6t
xi108 net561 net577 net550 sram_6t
xi107 bl2 bl2bar net550 sram_6t
xi106 net559 net575 net550 sram_6t
xi105 net572 net588 net550 sram_6t
xi96 net571 net587 net550 sram_6t
xi63 bl1 bl1bar net544 sram_6t
xi62 net569 net585 net544 sram_6t
xi61 net568 net584 net544 sram_6t
xi60 net652 net583 net544 sram_6t
xi59 bl0 bl0bar net544 sram_6t
xi58 net565 net581 net544 sram_6t
xi57 net558 net574 net544 sram_6t
xi56 bl1 bl1bar net546 sram_6t
xi13 net652 net583 net555 sram_6t
xi197 net557 net573 net548 sram_6t
xi192 net557 net573 net551 sram_6t
xi191 net557 net573 net555 sram_6t
xi190 net557 net573 net556 sram_6t
xi189 net557 net573 net655 sram_6t
xi40 bl1 bl1bar net548 sram_6t
xi39 net569 net585 net548 sram_6t
xi38 net568 net584 net548 sram_6t
xi37 net652 net583 net548 sram_6t
xi36 bl0 bl0bar net548 sram_6t
xi35 net565 net581 net548 sram_6t
xi34 net558 net574 net548 sram_6t
xi31 bl1 bl1bar net551 sram_6t
xi30 net569 net585 net551 sram_6t
xi29 net568 net584 net551 sram_6t
xi28 net652 net583 net551 sram_6t
xi27 bl0 bl0bar net551 sram_6t
xi26 net565 net581 net551 sram_6t
xi25 net558 net574 net551 sram_6t
xi23 bl1 bl1bar net556 sram_6t
xi22 net569 net585 net556 sram_6t
xi21 net568 net584 net556 sram_6t
xi20 net652 net583 net556 sram_6t
xi19 bl0 bl0bar net556 sram_6t
xi18 net565 net581 net556 sram_6t
xi17 net558 net574 net556 sram_6t
xi16 bl1 bl1bar net555 sram_6t
xi15 net569 net585 net555 sram_6t
xi14 net568 net584 net555 sram_6t
xi12 bl0 bl0bar net555 sram_6t
xi11 net565 net581 net555 sram_6t
xi118 net562 net578 net546 sram_6t
xi10 net558 net574 net555 sram_6t
xi119 net563 net579 net546 sram_6t
xi120 bl3 bl3bar net546 sram_6t
xi121 net572 net588 net544 sram_6t
xi122 net559 net575 net544 sram_6t
xi123 bl2 bl2bar net544 sram_6t
xi7 bl1 bl1bar net655 sram_6t
xi124 net561 net577 net544 sram_6t
xi125 net562 net578 net544 sram_6t
xi126 net563 net579 net544 sram_6t
xi127 bl3 bl3bar net544 sram_6t
xi6 net569 net585 net655 sram_6t
xi5 net568 net584 net655 sram_6t
xi4 net652 net583 net655 sram_6t
xi193 net557 net573 net550 sram_6t
xi3 bl0 bl0bar net655 sram_6t
xi2 net565 net581 net655 sram_6t
xi1 net558 net574 net655 sram_6t
xi41 net558 net574 net550 sram_6t
xi42 net565 net581 net550 sram_6t
xi43 bl0 bl0bar net550 sram_6t
xi44 net652 net583 net550 sram_6t
xi45 net568 net584 net550 sram_6t
xi46 net569 net585 net550 sram_6t
xi198 net557 net573 net544 sram_6t
xi202 a<2> a<3> a<4> wlref net544 net546 net550 net548 net551 net556 net555
+ net655 static_row_decoder_3by8
xi204 net557 net573 net558 net574 net565 net581 bl0 bl0bar net652 bl0 net568
+ net584 net569 net585 bl1 bl1bar net571 net587 net572 net588 net559 net575 bl2
+ bl2bar net561 net577 net562 net578 net563 net579 bl3 bl3bar net478 net476
+ net481 net479 2_driver 2_driverbar net487 net485 net490 net488 net493 net491
+ net496 net494 net499 net497 rs0 rs0bar rs1 rs1bar ws0 ws0bar ws1 ws1bar
+ columndecoder
xi206 d<1> net479 net481 write_driver
xi208 d<3> net485 net487 write_driver
xi205 d<0> net476 net478 write_driver
xi207 d<2> 2_driverbar 2_driver write_driver
xi211 net496 net494 read_dff2 read_circuit
xi212 net499 net497 read_dff3 read_circuit
xi209 net490 net488 read_dff0 read_circuit
xi210 net493 net491 read_dff1 read_circuit
xi215 read_dff3 q<3> net511 tspc_pos_ff
xi213 read_dff1 q<1> net511 tspc_pos_ff
xi214 read_dff2 q<2> net511 tspc_pos_ff
xi216 read_dff0 q<0> net511 tspc_pos_ff
xi217 a<0> a<1> net631 net613 net616 net619 wenb net622 net625 net628 net634
+ agen_unit
xi218 clk pc net659 wlref net511 wlref_pc
xi232 clk net622 net644 nand
xi233 clk net625 net646 nand
xi234 clk net628 net648 nand
xi236 clk net634 net650 nand
xi237 net636 rs0 inv_highdrive
xi238 net638 rs0bar inv_highdrive
xi239 net640 rs1 inv_highdrive
xi240 net642 rs1bar inv_highdrive
xi241 net644 ws0 inv_highdrive
xi242 net646 ws0bar inv_highdrive
xi243 net648 ws1 inv_highdrive
xi244 net650 ws1bar inv_highdrive
xi229 net659 net613 net638 nor
xi230 net659 net616 net640 nor
xi231 net659 net619 net642 nor
xi235 net659 net631 net636 nor
.ends memory_array

********************************************************************************
* Library          : group8
* Cell             : tb2025_2_tree_decoder
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
c1 q<1> gnd! c=1f
c3 q<3> gnd! c=1f
c2 q<2> gnd! c=1f
c0 q<0> gnd! c=1f
r33 i_a<4> gnd! r=1meg
rdwenb i_wenb gnd! r=1meg
rdar1 i_a<3> gnd! r=1meg
rdar0 i_a<2> gnd! r=1meg
rdaw1 i_a<1> gnd! r=1meg
rdaw0 i_a<0> gnd! r=1meg
rddw3 i_d<3> gnd! r=1meg
rddw2 i_d<2> gnd! r=1meg
rddw1 i_d<1> gnd! r=1meg
rddw0 i_d<0> gnd! r=1meg
xi34 a<4> i_a<4> inputbuf
xi25 clk net35 inputbuf
xbwenb wenb i_wenb inputbuf
xbar1 a<3> i_a<3> inputbuf
xbar0 a<2> i_a<2> inputbuf
xbaw1 a<1> i_a<1> inputbuf
xbaw0 a<0> i_a<0> inputbuf
xbdw3 d<3> i_d<3> inputbuf
xbdw2 d<2> i_d<2> inputbuf
xbdw1 d<1> i_d<1> inputbuf
xbdw0 d<0> i_d<0> inputbuf
vclk net35 gnd! dc=0 pulse ( 0 'vdd' 0 'clkrise' 'clkrise' '(clkperiod/2)-clkrise' 'clkperiod'
+  )
vdd vdd! gnd! dc='vdd'
xi35 a<0> a<1> a<2> a<3> a<4> clk d<0> d<1> d<2> d<3> q<0> q<1> q<2> q<3> wenb
+ memory_array









.tran 0.1p 6n start=0
.option opfile=1 split_dp=1
.option probe=1
.probe tran v(*) level=1
.probe tran v(a<0>) v(a<1>) v(a<2>) v(a<3>) v(a<4>) v(clk) v(d<0>) v(d<1>)
+ v(d<2>) v(d<3>) v(q<0>) v(q<1>) v(q<2>) v(q<3>) v(wenb)








.end
