* PEX netlist file	Thu Apr 17 14:24:02 2025	Cmux2
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 1
.subckt nor 2 3 4 5 6 7 8 9 10
.ends nor
.subckt inv 2 3 4 5 6 7 8 9
.ends inv
.subckt nand 2 3 4 5 6 7 9 11 12 13
*.floating_nets 8 10 14 15
MM1 3 6 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=808 $Y=543  $PIN_XY=838,608,808,543,778,608 $DEVICE_ID=1003
MM2 4 5 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=640 $Y=522  $PIN_XY=670,608,640,522,610,608 $DEVICE_ID=1003
.ends nand
.subckt 2to4_decoder_static_filler_17 2 3 4 5 6 7 8 9
.ends 2to4_decoder_static_filler_17

* Hierarchy Level 0

* Top of hierarchy  cell=Cmux2
.subckt Cmux2 GND! VDD! BL0 IN0 OP0 IN0BAR OP0BAR BL1 BL2 BL3 12
+	RS1 14 RS1BAR 16 WS1BAR WS1 19 20 21 22 23
+	24 WS0BAR RS0BAR 27 RS0 WS0 30 31 32 33 34
+	35 36 37 BL0_BAR BL1_BAR BL2_BAR BL3_BAR 46 47 48 49
+	50 51 52 53 54 55 56 57 58 59 60
+	61 62 63 64 65 66 67 68 69 70 71
+	72 73 74 75 76 77
*.floating_nets 87
MM1 IN0BAR 24 BL3_BAR nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2574 $Y=2243  $PIN_XY=2604,2226,2574,2243,2544,2226 $DEVICE_ID=1001
MM2 35 WS0 108 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=273  $PIN_XY=2436,378,2406,273,2376,378 $DEVICE_ID=1001
MM3 IN0 24 BL3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2238 $Y=2243  $PIN_XY=2268,2226,2238,2243,2208,2226 $DEVICE_ID=1001
MM4 24 35 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2238 $Y=756  $PIN_XY=2268,672,2238,756,2208,672 $DEVICE_ID=1001
MM5 108 WS1 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=294  $PIN_XY=2268,378,2238,294,2208,378 $DEVICE_ID=1001
MM6 IN0BAR 23 BL2_BAR nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1902 $Y=2243  $PIN_XY=1932,2226,1902,2243,1872,2226 $DEVICE_ID=1001
MM7 33 WS1 107 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=273  $PIN_XY=1764,378,1734,273,1704,378 $DEVICE_ID=1001
MM8 IN0 23 BL2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1566 $Y=2243  $PIN_XY=1596,2226,1566,2243,1536,2226 $DEVICE_ID=1001
MM9 23 33 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1566 $Y=756  $PIN_XY=1596,672,1566,756,1536,672 $DEVICE_ID=1001
MM10 107 WS0BAR GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=294  $PIN_XY=1596,378,1566,294,1536,378 $DEVICE_ID=1001
MM11 IN0BAR 21 BL1_BAR nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1230 $Y=2243  $PIN_XY=1260,2226,1230,2243,1200,2226 $DEVICE_ID=1001
MM12 30 WS0 106 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=273  $PIN_XY=1092,378,1062,273,1032,378 $DEVICE_ID=1001
MM13 IN0 21 BL1 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=894 $Y=2243  $PIN_XY=924,2226,894,2243,864,2226 $DEVICE_ID=1001
MM14 21 30 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=894 $Y=756  $PIN_XY=924,672,894,756,864,672 $DEVICE_ID=1001
MM15 106 WS1BAR GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=294  $PIN_XY=924,378,894,294,864,378 $DEVICE_ID=1001
MM16 IN0BAR 19 BL0_BAR nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=558 $Y=2243  $PIN_XY=588,2226,558,2243,528,2226 $DEVICE_ID=1001
MM17 27 WS1BAR 105 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=273  $PIN_XY=420,378,390,273,360,378 $DEVICE_ID=1001
MM18 IN0 19 BL0 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=2243  $PIN_XY=252,2226,222,2243,192,2226 $DEVICE_ID=1001
MM19 19 27 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=756  $PIN_XY=252,672,222,756,192,672 $DEVICE_ID=1001
MM20 105 WS0BAR GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=294  $PIN_XY=252,378,222,294,192,378 $DEVICE_ID=1001
MM21 OP0BAR 37 BL3_BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2574 $Y=3628  $PIN_XY=2604,3614,2574,3628,2544,3614 $DEVICE_ID=1003
MM22 VDD! 12 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=1781  $PIN_XY=2436,1766,2406,1781,2376,1766 $DEVICE_ID=1003
MM23 12 RS1 112 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=1197  $PIN_XY=2436,1132,2406,1197,2376,1132 $DEVICE_ID=1003
MM24 VDD! 35 24 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2406 $Y=857  $PIN_XY=2436,842,2406,857,2376,842 $DEVICE_ID=1003
MM25 OP0 37 BL3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2238 $Y=3628  $PIN_XY=2268,3614,2238,3628,2208,3614 $DEVICE_ID=1003
MM26 34 12 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=1680  $PIN_XY=2268,1766,2238,1680,2208,1766 $DEVICE_ID=1003
MM27 112 RS0 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=1218  $PIN_XY=2268,1132,2238,1218,2208,1132 $DEVICE_ID=1003
MM28 24 35 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2238 $Y=756  $PIN_XY=2268,842,2238,756,2208,842 $DEVICE_ID=1003
MM29 OP0BAR 36 BL2_BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1902 $Y=3628  $PIN_XY=1932,3614,1902,3628,1872,3614 $DEVICE_ID=1003
MM30 VDD! 31 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=1781  $PIN_XY=1764,1766,1734,1781,1704,1766 $DEVICE_ID=1003
MM31 31 RS1 111 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=1197  $PIN_XY=1764,1132,1734,1197,1704,1132 $DEVICE_ID=1003
MM32 VDD! 33 23 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1734 $Y=857  $PIN_XY=1764,842,1734,857,1704,842 $DEVICE_ID=1003
MM33 OP0 36 BL2 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1566 $Y=3628  $PIN_XY=1596,3614,1566,3628,1536,3614 $DEVICE_ID=1003
MM34 32 31 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=1680  $PIN_XY=1596,1766,1566,1680,1536,1766 $DEVICE_ID=1003
MM35 111 RS0BAR VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=1218  $PIN_XY=1596,1132,1566,1218,1536,1132 $DEVICE_ID=1003
MM36 23 33 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1566 $Y=756  $PIN_XY=1596,842,1566,756,1536,842 $DEVICE_ID=1003
MM37 OP0BAR 22 BL1_BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1230 $Y=3628  $PIN_XY=1260,3614,1230,3628,1200,3614 $DEVICE_ID=1003
MM38 VDD! 14 22 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=1781  $PIN_XY=1092,1766,1062,1781,1032,1766 $DEVICE_ID=1003
MM39 14 RS1BAR 110 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=1197  $PIN_XY=1092,1132,1062,1197,1032,1132 $DEVICE_ID=1003
MM40 VDD! 30 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1062 $Y=857  $PIN_XY=1092,842,1062,857,1032,842 $DEVICE_ID=1003
MM41 OP0 22 BL1 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=894 $Y=3628  $PIN_XY=924,3614,894,3628,864,3614 $DEVICE_ID=1003
MM42 22 14 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=1680  $PIN_XY=924,1766,894,1680,864,1766 $DEVICE_ID=1003
MM43 110 RS0 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=1218  $PIN_XY=924,1132,894,1218,864,1132 $DEVICE_ID=1003
MM44 21 30 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=894 $Y=756  $PIN_XY=924,842,894,756,864,842 $DEVICE_ID=1003
MM45 OP0BAR 20 BL0_BAR pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=558 $Y=3628  $PIN_XY=588,3614,558,3628,528,3614 $DEVICE_ID=1003
MM46 VDD! 16 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=1781  $PIN_XY=420,1766,390,1781,360,1766 $DEVICE_ID=1003
MM47 16 RS1BAR 109 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=1197  $PIN_XY=420,1132,390,1197,360,1132 $DEVICE_ID=1003
MM48 VDD! 27 19 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=857  $PIN_XY=420,842,390,857,360,842 $DEVICE_ID=1003
MM49 OP0 20 BL0 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=3628  $PIN_XY=252,3614,222,3628,192,3614 $DEVICE_ID=1003
MM50 20 16 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=1680  $PIN_XY=252,1766,222,1680,192,1766 $DEVICE_ID=1003
MM51 109 RS0BAR VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=1218  $PIN_XY=252,1132,222,1218,192,1132 $DEVICE_ID=1003
MM52 19 27 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=756  $PIN_XY=252,842,222,756,192,842 $DEVICE_ID=1003
XXA327B7031 GND! VDD! 32 31 RS0BAR 44 GND! 89 inv $T=1344 1386 0 0 $X=1344 $Y=1386
XXA327B7032 GND! VDD! 34 12 RS0 45 GND! 90 inv $T=2016 1386 0 0 $X=2016 $Y=1386
XXA327B7033 GND! VDD! 22 14 RS0 43 GND! 91 inv $T=672 1386 0 0 $X=672 $Y=1386
XXA327B7034 GND! VDD! 20 16 RS0BAR 42 GND! 92 inv $T=0 1386 0 0 $X=0 $Y=1386
XXA327B7035 GND! VDD! 24 35 WS1 81 GND! 93 inv $T=2016 462 0 0 $X=2016 $Y=462
XXA327B7036 GND! VDD! 23 33 WS0BAR 80 GND! 94 inv $T=1344 462 0 0 $X=1344 $Y=462
XXA327B7037 GND! VDD! 21 30 WS1BAR 79 GND! 95 inv $T=672 462 0 0 $X=672 $Y=462
XXA327B7038 GND! VDD! 19 27 WS0BAR 78 GND! 96 inv $T=0 462 0 0 $X=0 $Y=462
XXA327B7039 GND! VDD! 97 VDD! GND! _GENERATED_113 82 88 2to4_decoder_static_filler_17 $T=3132 588 0 180 $X=2688 $Y=-2
XXA327B70310 GND! VDD! GND! _GENERATED_114 98 VDD! 82 GND! 2to4_decoder_static_filler_17 $T=2688 462 0 0 $X=2688 $Y=462
XXA327B70311 GND! VDD! 99 VDD! GND! _GENERATED_115 83 GND! 2to4_decoder_static_filler_17 $T=3132 1512 0 180 $X=2688 $Y=922
XXA327B70312 GND! VDD! GND! _GENERATED_116 100 VDD! 83 GND! 2to4_decoder_static_filler_17 $T=2688 1386 0 0 $X=2688 $Y=1386
XXA327B70313 GND! VDD! 101 VDD! GND! _GENERATED_117 84 GND! 2to4_decoder_static_filler_17 $T=3132 2436 0 180 $X=2688 $Y=1846
XXA327B70314 GND! VDD! GND! _GENERATED_118 102 VDD! 84 BL0 2to4_decoder_static_filler_17 $T=2688 2310 0 0 $X=2688 $Y=2310
XXA327B70315 GND! VDD! 103 VDD! GND! _GENERATED_119 85 BL0 2to4_decoder_static_filler_17 $T=3132 3360 0 180 $X=2688 $Y=2770
XXA327B70316 GND! VDD! GND! _GENERATED_120 104 VDD! 85 OP0 2to4_decoder_static_filler_17 $T=2688 3234 0 0 $X=2688 $Y=3234
XXA327B70317 GND! VDD! 12 RS1 RS0 12 35 35 112 nor $T=1388 1514 1 0 $X=2016 $Y=922
XXA327B70318 GND! VDD! 31 RS1 RS0BAR 31 33 33 111 nor $T=716 1514 1 0 $X=1343 $Y=922
XXA327B70319 GND! VDD! 14 RS1BAR RS0 14 30 30 110 nor $T=44 1514 1 0 $X=672 $Y=922
XXA327B70320 GND! VDD! 16 RS1BAR RS0BAR 16 27 27 109 nor $T=-628 1514 1 0 $X=0 $Y=922
XXA327B70321 GND! VDD! 27 WS0BAR WS1BAR 27 105 82 86 88 nand $T=-418 816 1 0 $X=0 $Y=-2
XXA327B70322 GND! VDD! 30 WS1BAR WS0 30 106 82 86 88 nand $T=254 816 1 0 $X=671 $Y=-2
XXA327B70323 GND! VDD! 33 WS0BAR WS1 33 107 82 86 88 nand $T=926 816 1 0 $X=1344 $Y=-2
XXA327B70324 GND! VDD! 35 WS1 WS0 35 108 82 86 88 nand $T=1598 816 1 0 $X=2016 $Y=-2
.ends Cmux2
