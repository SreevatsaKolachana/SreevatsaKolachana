* PEX netlist file	Sat Apr 12 15:24:33 2025	memory_array_8by16
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 1
.subckt sram_6t 2 3 4 5 6 7 8 9 10 11 12
+	13 16 17 18
*.floating_nets 14 15 19 20
MM1 3 6 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=366 $Y=756  $PIN_XY=396,670,366,756,336,670 $DEVICE_ID=1003
MM2 6 7 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=198 $Y=294  $PIN_XY=228,380,198,294,168,380 $DEVICE_ID=1003
.ends sram_6t
.subckt sram_filler 2 3 4 5
.ends sram_filler

* Hierarchy Level 0

* Top of hierarchy  cell=memory_array_8by16
.subckt memory_array_8by16 GND! VDD! WL<0> WL<1> WL<2> WL<3> WL<4> WL<5> WL<6> WL<7> BLB<1>
+	BL<1> BLB<0> BL<0> BLB<4> BL<4> BLB<2> BL<2> BLB<3> BL<3> BLB<5> BL<5>
+	BLB<7> BL<7> BLB<6> BL<6> BLB<8> BL<8> BLB<9> BL<9> BLB<10> BL<10> BLB<11>
+	BL<11> BLB<12> BL<12> BLB<14> BL<14> BLB<15> BL<15> BLB<13> BL<13>
MM1 GND! 368 264 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=7242  $PIN_XY=9076,7326,9046,7242,9016,7326 $DEVICE_ID=1001
MM2 BL<15> WL<7> 368 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=6693  $PIN_XY=9076,6696,9046,6693,9016,6696 $DEVICE_ID=1001
MM3 GND! 265 254 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=6318  $PIN_XY=9076,6402,9046,6318,9016,6402 $DEVICE_ID=1001
MM4 BL<15> WL<6> 265 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=5769  $PIN_XY=9076,5772,9046,5769,9016,5772 $DEVICE_ID=1001
MM5 GND! 255 248 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=5394  $PIN_XY=9076,5478,9046,5394,9016,5478 $DEVICE_ID=1001
MM6 BL<15> WL<5> 255 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=4845  $PIN_XY=9076,4848,9046,4845,9016,4848 $DEVICE_ID=1001
MM7 GND! 249 158 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=4470  $PIN_XY=9076,4554,9046,4470,9016,4554 $DEVICE_ID=1001
MM8 264 WL<7> BLB<15> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=7329  $PIN_XY=8908,7326,8878,7329,8848,7326 $DEVICE_ID=1001
MM9 368 264 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=6780  $PIN_XY=8908,6696,8878,6780,8848,6696 $DEVICE_ID=1001
MM10 254 WL<6> BLB<15> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=6405  $PIN_XY=8908,6402,8878,6405,8848,6402 $DEVICE_ID=1001
MM11 265 254 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=5856  $PIN_XY=8908,5772,8878,5856,8848,5772 $DEVICE_ID=1001
MM12 248 WL<5> BLB<15> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=5481  $PIN_XY=8908,5478,8878,5481,8848,5478 $DEVICE_ID=1001
MM13 255 248 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=4932  $PIN_XY=8908,4848,8878,4932,8848,4848 $DEVICE_ID=1001
MM14 158 WL<4> BLB<15> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=4557  $PIN_XY=8908,4554,8878,4557,8848,4554 $DEVICE_ID=1001
MM15 GND! 371 266 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=7242  $PIN_XY=8572,7326,8542,7242,8512,7326 $DEVICE_ID=1001
MM16 BL<14> WL<7> 371 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=6693  $PIN_XY=8572,6696,8542,6693,8512,6696 $DEVICE_ID=1001
MM17 GND! 267 252 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=6318  $PIN_XY=8572,6402,8542,6318,8512,6402 $DEVICE_ID=1001
MM18 BL<14> WL<6> 267 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=5769  $PIN_XY=8572,5772,8542,5769,8512,5772 $DEVICE_ID=1001
MM19 GND! 253 250 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=5394  $PIN_XY=8572,5478,8542,5394,8512,5478 $DEVICE_ID=1001
MM20 BL<14> WL<5> 253 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=4845  $PIN_XY=8572,4848,8542,4845,8512,4848 $DEVICE_ID=1001
MM21 GND! 251 156 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=4470  $PIN_XY=8572,4554,8542,4470,8512,4554 $DEVICE_ID=1001
MM22 266 WL<7> BLB<14> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=7329  $PIN_XY=8404,7326,8374,7329,8344,7326 $DEVICE_ID=1001
MM23 371 266 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=6780  $PIN_XY=8404,6696,8374,6780,8344,6696 $DEVICE_ID=1001
MM24 252 WL<6> BLB<14> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=6405  $PIN_XY=8404,6402,8374,6405,8344,6402 $DEVICE_ID=1001
MM25 267 252 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=5856  $PIN_XY=8404,5772,8374,5856,8344,5772 $DEVICE_ID=1001
MM26 250 WL<5> BLB<14> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=5481  $PIN_XY=8404,5478,8374,5481,8344,5478 $DEVICE_ID=1001
MM27 253 250 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=4932  $PIN_XY=8404,4848,8374,4932,8344,4848 $DEVICE_ID=1001
MM28 156 WL<4> BLB<14> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=4557  $PIN_XY=8404,4554,8374,4557,8344,4554 $DEVICE_ID=1001
MM29 GND! 365 262 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=7242  $PIN_XY=8068,7326,8038,7242,8008,7326 $DEVICE_ID=1001
MM30 BL<13> WL<7> 365 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=6693  $PIN_XY=8068,6696,8038,6693,8008,6696 $DEVICE_ID=1001
MM31 GND! 263 256 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=6318  $PIN_XY=8068,6402,8038,6318,8008,6402 $DEVICE_ID=1001
MM32 BL<13> WL<6> 263 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=5769  $PIN_XY=8068,5772,8038,5769,8008,5772 $DEVICE_ID=1001
MM33 GND! 257 246 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=5394  $PIN_XY=8068,5478,8038,5394,8008,5478 $DEVICE_ID=1001
MM34 BL<13> WL<5> 257 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=4845  $PIN_XY=8068,4848,8038,4845,8008,4848 $DEVICE_ID=1001
MM35 GND! 247 160 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=4470  $PIN_XY=8068,4554,8038,4470,8008,4554 $DEVICE_ID=1001
MM36 262 WL<7> BLB<13> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=7329  $PIN_XY=7900,7326,7870,7329,7840,7326 $DEVICE_ID=1001
MM37 365 262 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=6780  $PIN_XY=7900,6696,7870,6780,7840,6696 $DEVICE_ID=1001
MM38 256 WL<6> BLB<13> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=6405  $PIN_XY=7900,6402,7870,6405,7840,6402 $DEVICE_ID=1001
MM39 263 256 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=5856  $PIN_XY=7900,5772,7870,5856,7840,5772 $DEVICE_ID=1001
MM40 246 WL<5> BLB<13> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=5481  $PIN_XY=7900,5478,7870,5481,7840,5478 $DEVICE_ID=1001
MM41 257 246 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=4932  $PIN_XY=7900,4848,7870,4932,7840,4848 $DEVICE_ID=1001
MM42 160 WL<4> BLB<13> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=4557  $PIN_XY=7900,4554,7870,4557,7840,4554 $DEVICE_ID=1001
MM43 GND! 362 260 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=7242  $PIN_XY=7564,7326,7534,7242,7504,7326 $DEVICE_ID=1001
MM44 BL<12> WL<7> 362 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=6693  $PIN_XY=7564,6696,7534,6693,7504,6696 $DEVICE_ID=1001
MM45 GND! 261 258 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=6318  $PIN_XY=7564,6402,7534,6318,7504,6402 $DEVICE_ID=1001
MM46 BL<12> WL<6> 261 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=5769  $PIN_XY=7564,5772,7534,5769,7504,5772 $DEVICE_ID=1001
MM47 GND! 259 244 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=5394  $PIN_XY=7564,5478,7534,5394,7504,5478 $DEVICE_ID=1001
MM48 BL<12> WL<5> 259 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=4845  $PIN_XY=7564,4848,7534,4845,7504,4848 $DEVICE_ID=1001
MM49 GND! 245 162 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=4470  $PIN_XY=7564,4554,7534,4470,7504,4554 $DEVICE_ID=1001
MM50 260 WL<7> BLB<12> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=7329  $PIN_XY=7396,7326,7366,7329,7336,7326 $DEVICE_ID=1001
MM51 362 260 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=6780  $PIN_XY=7396,6696,7366,6780,7336,6696 $DEVICE_ID=1001
MM52 258 WL<6> BLB<12> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=6405  $PIN_XY=7396,6402,7366,6405,7336,6402 $DEVICE_ID=1001
MM53 261 258 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=5856  $PIN_XY=7396,5772,7366,5856,7336,5772 $DEVICE_ID=1001
MM54 244 WL<5> BLB<12> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=5481  $PIN_XY=7396,5478,7366,5481,7336,5478 $DEVICE_ID=1001
MM55 259 244 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=4932  $PIN_XY=7396,4848,7366,4932,7336,4848 $DEVICE_ID=1001
MM56 162 WL<4> BLB<12> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=4557  $PIN_XY=7396,4554,7366,4557,7336,4554 $DEVICE_ID=1001
MM57 GND! 356 240 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=7242  $PIN_XY=6724,7326,6694,7242,6664,7326 $DEVICE_ID=1001
MM58 BL<11> WL<7> 356 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=6693  $PIN_XY=6724,6696,6694,6693,6664,6696 $DEVICE_ID=1001
MM59 GND! 241 234 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=6318  $PIN_XY=6724,6402,6694,6318,6664,6402 $DEVICE_ID=1001
MM60 BL<11> WL<6> 241 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=5769  $PIN_XY=6724,5772,6694,5769,6664,5772 $DEVICE_ID=1001
MM61 GND! 235 228 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=5394  $PIN_XY=6724,5478,6694,5394,6664,5478 $DEVICE_ID=1001
MM62 BL<11> WL<5> 235 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=4845  $PIN_XY=6724,4848,6694,4845,6664,4848 $DEVICE_ID=1001
MM63 GND! 229 130 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=4470  $PIN_XY=6724,4554,6694,4470,6664,4554 $DEVICE_ID=1001
MM64 240 WL<7> BLB<11> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=7329  $PIN_XY=6556,7326,6526,7329,6496,7326 $DEVICE_ID=1001
MM65 356 240 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=6780  $PIN_XY=6556,6696,6526,6780,6496,6696 $DEVICE_ID=1001
MM66 234 WL<6> BLB<11> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=6405  $PIN_XY=6556,6402,6526,6405,6496,6402 $DEVICE_ID=1001
MM67 241 234 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=5856  $PIN_XY=6556,5772,6526,5856,6496,5772 $DEVICE_ID=1001
MM68 228 WL<5> BLB<11> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=5481  $PIN_XY=6556,5478,6526,5481,6496,5478 $DEVICE_ID=1001
MM69 235 228 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=4932  $PIN_XY=6556,4848,6526,4932,6496,4848 $DEVICE_ID=1001
MM70 130 WL<4> BLB<11> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=4557  $PIN_XY=6556,4554,6526,4557,6496,4554 $DEVICE_ID=1001
MM71 GND! 353 238 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=7242  $PIN_XY=6220,7326,6190,7242,6160,7326 $DEVICE_ID=1001
MM72 BL<10> WL<7> 353 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=6693  $PIN_XY=6220,6696,6190,6693,6160,6696 $DEVICE_ID=1001
MM73 GND! 239 236 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=6318  $PIN_XY=6220,6402,6190,6318,6160,6402 $DEVICE_ID=1001
MM74 BL<10> WL<6> 239 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=5769  $PIN_XY=6220,5772,6190,5769,6160,5772 $DEVICE_ID=1001
MM75 GND! 237 226 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=5394  $PIN_XY=6220,5478,6190,5394,6160,5478 $DEVICE_ID=1001
MM76 BL<10> WL<5> 237 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=4845  $PIN_XY=6220,4848,6190,4845,6160,4848 $DEVICE_ID=1001
MM77 GND! 227 132 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=4470  $PIN_XY=6220,4554,6190,4470,6160,4554 $DEVICE_ID=1001
MM78 238 WL<7> BLB<10> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=7329  $PIN_XY=6052,7326,6022,7329,5992,7326 $DEVICE_ID=1001
MM79 353 238 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=6780  $PIN_XY=6052,6696,6022,6780,5992,6696 $DEVICE_ID=1001
MM80 236 WL<6> BLB<10> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=6405  $PIN_XY=6052,6402,6022,6405,5992,6402 $DEVICE_ID=1001
MM81 239 236 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=5856  $PIN_XY=6052,5772,6022,5856,5992,5772 $DEVICE_ID=1001
MM82 226 WL<5> BLB<10> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=5481  $PIN_XY=6052,5478,6022,5481,5992,5478 $DEVICE_ID=1001
MM83 237 226 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=4932  $PIN_XY=6052,4848,6022,4932,5992,4848 $DEVICE_ID=1001
MM84 132 WL<4> BLB<10> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=4557  $PIN_XY=6052,4554,6022,4557,5992,4554 $DEVICE_ID=1001
MM85 GND! 359 242 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=7242  $PIN_XY=5716,7326,5686,7242,5656,7326 $DEVICE_ID=1001
MM86 BL<9> WL<7> 359 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=6693  $PIN_XY=5716,6696,5686,6693,5656,6696 $DEVICE_ID=1001
MM87 GND! 243 232 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=6318  $PIN_XY=5716,6402,5686,6318,5656,6402 $DEVICE_ID=1001
MM88 BL<9> WL<6> 243 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=5769  $PIN_XY=5716,5772,5686,5769,5656,5772 $DEVICE_ID=1001
MM89 GND! 233 230 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=5394  $PIN_XY=5716,5478,5686,5394,5656,5478 $DEVICE_ID=1001
MM90 BL<9> WL<5> 233 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=4845  $PIN_XY=5716,4848,5686,4845,5656,4848 $DEVICE_ID=1001
MM91 GND! 231 128 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=4470  $PIN_XY=5716,4554,5686,4470,5656,4554 $DEVICE_ID=1001
MM92 242 WL<7> BLB<9> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=7329  $PIN_XY=5548,7326,5518,7329,5488,7326 $DEVICE_ID=1001
MM93 359 242 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=6780  $PIN_XY=5548,6696,5518,6780,5488,6696 $DEVICE_ID=1001
MM94 232 WL<6> BLB<9> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=6405  $PIN_XY=5548,6402,5518,6405,5488,6402 $DEVICE_ID=1001
MM95 243 232 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=5856  $PIN_XY=5548,5772,5518,5856,5488,5772 $DEVICE_ID=1001
MM96 230 WL<5> BLB<9> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=5481  $PIN_XY=5548,5478,5518,5481,5488,5478 $DEVICE_ID=1001
MM97 233 230 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=4932  $PIN_XY=5548,4848,5518,4932,5488,4848 $DEVICE_ID=1001
MM98 128 WL<4> BLB<9> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=4557  $PIN_XY=5548,4554,5518,4557,5488,4554 $DEVICE_ID=1001
MM99 GND! 350 224 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=7242  $PIN_XY=5212,7326,5182,7242,5152,7326 $DEVICE_ID=1001
MM100 BL<8> WL<7> 350 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=6693  $PIN_XY=5212,6696,5182,6693,5152,6696 $DEVICE_ID=1001
MM101 GND! 225 214 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=6318  $PIN_XY=5212,6402,5182,6318,5152,6402 $DEVICE_ID=1001
MM102 BL<8> WL<6> 225 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=5769  $PIN_XY=5212,5772,5182,5769,5152,5772 $DEVICE_ID=1001
MM103 GND! 215 212 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=5394  $PIN_XY=5212,5478,5182,5394,5152,5478 $DEVICE_ID=1001
MM104 BL<8> WL<5> 215 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=4845  $PIN_XY=5212,4848,5182,4845,5152,4848 $DEVICE_ID=1001
MM105 GND! 213 104 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=4470  $PIN_XY=5212,4554,5182,4470,5152,4554 $DEVICE_ID=1001
MM106 224 WL<7> BLB<8> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=7329  $PIN_XY=5044,7326,5014,7329,4984,7326 $DEVICE_ID=1001
MM107 350 224 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=6780  $PIN_XY=5044,6696,5014,6780,4984,6696 $DEVICE_ID=1001
MM108 214 WL<6> BLB<8> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=6405  $PIN_XY=5044,6402,5014,6405,4984,6402 $DEVICE_ID=1001
MM109 225 214 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=5856  $PIN_XY=5044,5772,5014,5856,4984,5772 $DEVICE_ID=1001
MM110 212 WL<5> BLB<8> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=5481  $PIN_XY=5044,5478,5014,5481,4984,5478 $DEVICE_ID=1001
MM111 215 212 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=4932  $PIN_XY=5044,4848,5014,4932,4984,4848 $DEVICE_ID=1001
MM112 104 WL<4> BLB<8> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=4557  $PIN_XY=5044,4554,5014,4557,4984,4554 $DEVICE_ID=1001
MM113 GND! 347 222 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=7242  $PIN_XY=4372,7326,4342,7242,4312,7326 $DEVICE_ID=1001
MM114 BL<7> WL<7> 347 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=6693  $PIN_XY=4372,6696,4342,6693,4312,6696 $DEVICE_ID=1001
MM115 GND! 223 216 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=6318  $PIN_XY=4372,6402,4342,6318,4312,6402 $DEVICE_ID=1001
MM116 BL<7> WL<6> 223 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=5769  $PIN_XY=4372,5772,4342,5769,4312,5772 $DEVICE_ID=1001
MM117 GND! 217 210 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=5394  $PIN_XY=4372,5478,4342,5394,4312,5478 $DEVICE_ID=1001
MM118 BL<7> WL<5> 217 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=4845  $PIN_XY=4372,4848,4342,4845,4312,4848 $DEVICE_ID=1001
MM119 GND! 211 106 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=4470  $PIN_XY=4372,4554,4342,4470,4312,4554 $DEVICE_ID=1001
MM120 222 WL<7> BLB<7> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=7329  $PIN_XY=4204,7326,4174,7329,4144,7326 $DEVICE_ID=1001
MM121 347 222 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=6780  $PIN_XY=4204,6696,4174,6780,4144,6696 $DEVICE_ID=1001
MM122 216 WL<6> BLB<7> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=6405  $PIN_XY=4204,6402,4174,6405,4144,6402 $DEVICE_ID=1001
MM123 223 216 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=5856  $PIN_XY=4204,5772,4174,5856,4144,5772 $DEVICE_ID=1001
MM124 210 WL<5> BLB<7> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=5481  $PIN_XY=4204,5478,4174,5481,4144,5478 $DEVICE_ID=1001
MM125 217 210 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=4932  $PIN_XY=4204,4848,4174,4932,4144,4848 $DEVICE_ID=1001
MM126 106 WL<4> BLB<7> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=4557  $PIN_XY=4204,4554,4174,4557,4144,4554 $DEVICE_ID=1001
MM127 GND! 344 220 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=7242  $PIN_XY=3868,7326,3838,7242,3808,7326 $DEVICE_ID=1001
MM128 BL<6> WL<7> 344 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=6693  $PIN_XY=3868,6696,3838,6693,3808,6696 $DEVICE_ID=1001
MM129 GND! 221 218 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=6318  $PIN_XY=3868,6402,3838,6318,3808,6402 $DEVICE_ID=1001
MM130 BL<6> WL<6> 221 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=5769  $PIN_XY=3868,5772,3838,5769,3808,5772 $DEVICE_ID=1001
MM131 GND! 219 208 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=5394  $PIN_XY=3868,5478,3838,5394,3808,5478 $DEVICE_ID=1001
MM132 BL<6> WL<5> 219 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=4845  $PIN_XY=3868,4848,3838,4845,3808,4848 $DEVICE_ID=1001
MM133 GND! 209 108 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=4470  $PIN_XY=3868,4554,3838,4470,3808,4554 $DEVICE_ID=1001
MM134 220 WL<7> BLB<6> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=7329  $PIN_XY=3700,7326,3670,7329,3640,7326 $DEVICE_ID=1001
MM135 344 220 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=6780  $PIN_XY=3700,6696,3670,6780,3640,6696 $DEVICE_ID=1001
MM136 218 WL<6> BLB<6> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=6405  $PIN_XY=3700,6402,3670,6405,3640,6402 $DEVICE_ID=1001
MM137 221 218 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=5856  $PIN_XY=3700,5772,3670,5856,3640,5772 $DEVICE_ID=1001
MM138 208 WL<5> BLB<6> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=5481  $PIN_XY=3700,5478,3670,5481,3640,5478 $DEVICE_ID=1001
MM139 219 208 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=4932  $PIN_XY=3700,4848,3670,4932,3640,4848 $DEVICE_ID=1001
MM140 108 WL<4> BLB<6> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=4557  $PIN_XY=3700,4554,3670,4557,3640,4554 $DEVICE_ID=1001
MM141 GND! 338 204 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=7242  $PIN_XY=3364,7326,3334,7242,3304,7326 $DEVICE_ID=1001
MM142 BL<5> WL<7> 338 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=6693  $PIN_XY=3364,6696,3334,6693,3304,6696 $DEVICE_ID=1001
MM143 GND! 205 200 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=6318  $PIN_XY=3364,6402,3334,6318,3304,6402 $DEVICE_ID=1001
MM144 BL<5> WL<6> 205 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=5769  $PIN_XY=3364,5772,3334,5769,3304,5772 $DEVICE_ID=1001
MM145 GND! 201 192 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=5394  $PIN_XY=3364,5478,3334,5394,3304,5478 $DEVICE_ID=1001
MM146 BL<5> WL<5> 201 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=4845  $PIN_XY=3364,4848,3334,4845,3304,4848 $DEVICE_ID=1001
MM147 GND! 193 82 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=4470  $PIN_XY=3364,4554,3334,4470,3304,4554 $DEVICE_ID=1001
MM148 204 WL<7> BLB<5> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=7329  $PIN_XY=3196,7326,3166,7329,3136,7326 $DEVICE_ID=1001
MM149 338 204 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=6780  $PIN_XY=3196,6696,3166,6780,3136,6696 $DEVICE_ID=1001
MM150 200 WL<6> BLB<5> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=6405  $PIN_XY=3196,6402,3166,6405,3136,6402 $DEVICE_ID=1001
MM151 205 200 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=5856  $PIN_XY=3196,5772,3166,5856,3136,5772 $DEVICE_ID=1001
MM152 192 WL<5> BLB<5> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=5481  $PIN_XY=3196,5478,3166,5481,3136,5478 $DEVICE_ID=1001
MM153 201 192 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=4932  $PIN_XY=3196,4848,3166,4932,3136,4848 $DEVICE_ID=1001
MM154 82 WL<4> BLB<5> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=4557  $PIN_XY=3196,4554,3166,4557,3136,4554 $DEVICE_ID=1001
MM155 GND! 341 206 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=7242  $PIN_XY=2860,7326,2830,7242,2800,7326 $DEVICE_ID=1001
MM156 BL<4> WL<7> 341 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=6693  $PIN_XY=2860,6696,2830,6693,2800,6696 $DEVICE_ID=1001
MM157 GND! 207 198 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=6318  $PIN_XY=2860,6402,2830,6318,2800,6402 $DEVICE_ID=1001
MM158 BL<4> WL<6> 207 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=5769  $PIN_XY=2860,5772,2830,5769,2800,5772 $DEVICE_ID=1001
MM159 GND! 199 194 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=5394  $PIN_XY=2860,5478,2830,5394,2800,5478 $DEVICE_ID=1001
MM160 BL<4> WL<5> 199 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=4845  $PIN_XY=2860,4848,2830,4845,2800,4848 $DEVICE_ID=1001
MM161 GND! 195 80 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=4470  $PIN_XY=2860,4554,2830,4470,2800,4554 $DEVICE_ID=1001
MM162 206 WL<7> BLB<4> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=7329  $PIN_XY=2692,7326,2662,7329,2632,7326 $DEVICE_ID=1001
MM163 341 206 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=6780  $PIN_XY=2692,6696,2662,6780,2632,6696 $DEVICE_ID=1001
MM164 198 WL<6> BLB<4> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=6405  $PIN_XY=2692,6402,2662,6405,2632,6402 $DEVICE_ID=1001
MM165 207 198 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=5856  $PIN_XY=2692,5772,2662,5856,2632,5772 $DEVICE_ID=1001
MM166 194 WL<5> BLB<4> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=5481  $PIN_XY=2692,5478,2662,5481,2632,5478 $DEVICE_ID=1001
MM167 199 194 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=4932  $PIN_XY=2692,4848,2662,4932,2632,4848 $DEVICE_ID=1001
MM168 80 WL<4> BLB<4> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=4557  $PIN_XY=2692,4554,2662,4557,2632,4554 $DEVICE_ID=1001
MM169 GND! 335 196 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=7242  $PIN_XY=2020,7326,1990,7242,1960,7326 $DEVICE_ID=1001
MM170 BL<3> WL<7> 335 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=6693  $PIN_XY=2020,6696,1990,6693,1960,6696 $DEVICE_ID=1001
MM171 GND! 197 202 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=6318  $PIN_XY=2020,6402,1990,6318,1960,6402 $DEVICE_ID=1001
MM172 BL<3> WL<6> 197 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=5769  $PIN_XY=2020,5772,1990,5769,1960,5772 $DEVICE_ID=1001
MM173 GND! 203 190 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=5394  $PIN_XY=2020,5478,1990,5394,1960,5478 $DEVICE_ID=1001
MM174 BL<3> WL<5> 203 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=4845  $PIN_XY=2020,4848,1990,4845,1960,4848 $DEVICE_ID=1001
MM175 GND! 191 90 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=4470  $PIN_XY=2020,4554,1990,4470,1960,4554 $DEVICE_ID=1001
MM176 196 WL<7> BLB<3> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=7329  $PIN_XY=1852,7326,1822,7329,1792,7326 $DEVICE_ID=1001
MM177 335 196 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=6780  $PIN_XY=1852,6696,1822,6780,1792,6696 $DEVICE_ID=1001
MM178 202 WL<6> BLB<3> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=6405  $PIN_XY=1852,6402,1822,6405,1792,6402 $DEVICE_ID=1001
MM179 197 202 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=5856  $PIN_XY=1852,5772,1822,5856,1792,5772 $DEVICE_ID=1001
MM180 190 WL<5> BLB<3> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=5481  $PIN_XY=1852,5478,1822,5481,1792,5478 $DEVICE_ID=1001
MM181 203 190 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=4932  $PIN_XY=1852,4848,1822,4932,1792,4848 $DEVICE_ID=1001
MM182 90 WL<4> BLB<3> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=4557  $PIN_XY=1852,4554,1822,4557,1792,4554 $DEVICE_ID=1001
MM183 GND! 332 182 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=7242  $PIN_XY=1516,7326,1486,7242,1456,7326 $DEVICE_ID=1001
MM184 BL<2> WL<7> 332 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=6693  $PIN_XY=1516,6696,1486,6693,1456,6696 $DEVICE_ID=1001
MM185 GND! 183 184 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=6318  $PIN_XY=1516,6402,1486,6318,1456,6402 $DEVICE_ID=1001
MM186 BL<2> WL<6> 183 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=5769  $PIN_XY=1516,5772,1486,5769,1456,5772 $DEVICE_ID=1001
MM187 GND! 185 176 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=5394  $PIN_XY=1516,5478,1486,5394,1456,5478 $DEVICE_ID=1001
MM188 BL<2> WL<5> 185 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=4845  $PIN_XY=1516,4848,1486,4845,1456,4848 $DEVICE_ID=1001
MM189 GND! 177 62 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=4470  $PIN_XY=1516,4554,1486,4470,1456,4554 $DEVICE_ID=1001
MM190 182 WL<7> BLB<2> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=7329  $PIN_XY=1348,7326,1318,7329,1288,7326 $DEVICE_ID=1001
MM191 332 182 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=6780  $PIN_XY=1348,6696,1318,6780,1288,6696 $DEVICE_ID=1001
MM192 184 WL<6> BLB<2> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=6405  $PIN_XY=1348,6402,1318,6405,1288,6402 $DEVICE_ID=1001
MM193 183 184 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=5856  $PIN_XY=1348,5772,1318,5856,1288,5772 $DEVICE_ID=1001
MM194 176 WL<5> BLB<2> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=5481  $PIN_XY=1348,5478,1318,5481,1288,5478 $DEVICE_ID=1001
MM195 185 176 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=4932  $PIN_XY=1348,4848,1318,4932,1288,4848 $DEVICE_ID=1001
MM196 62 WL<4> BLB<2> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=4557  $PIN_XY=1348,4554,1318,4557,1288,4554 $DEVICE_ID=1001
MM197 GND! 329 180 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=7242  $PIN_XY=1012,7326,982,7242,952,7326 $DEVICE_ID=1001
MM198 BL<1> WL<7> 329 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=6693  $PIN_XY=1012,6696,982,6693,952,6696 $DEVICE_ID=1001
MM199 GND! 181 186 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=6318  $PIN_XY=1012,6402,982,6318,952,6402 $DEVICE_ID=1001
MM200 BL<1> WL<6> 181 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=5769  $PIN_XY=1012,5772,982,5769,952,5772 $DEVICE_ID=1001
MM201 GND! 187 174 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=5394  $PIN_XY=1012,5478,982,5394,952,5478 $DEVICE_ID=1001
MM202 BL<1> WL<5> 187 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=4845  $PIN_XY=1012,4848,982,4845,952,4848 $DEVICE_ID=1001
MM203 GND! 175 64 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=4470  $PIN_XY=1012,4554,982,4470,952,4554 $DEVICE_ID=1001
MM204 180 WL<7> BLB<1> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=7329  $PIN_XY=844,7326,814,7329,784,7326 $DEVICE_ID=1001
MM205 329 180 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=6780  $PIN_XY=844,6696,814,6780,784,6696 $DEVICE_ID=1001
MM206 186 WL<6> BLB<1> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=6405  $PIN_XY=844,6402,814,6405,784,6402 $DEVICE_ID=1001
MM207 181 186 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=5856  $PIN_XY=844,5772,814,5856,784,5772 $DEVICE_ID=1001
MM208 174 WL<5> BLB<1> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=5481  $PIN_XY=844,5478,814,5481,784,5478 $DEVICE_ID=1001
MM209 187 174 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=4932  $PIN_XY=844,4848,814,4932,784,4848 $DEVICE_ID=1001
MM210 64 WL<4> BLB<1> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=4557  $PIN_XY=844,4554,814,4557,784,4554 $DEVICE_ID=1001
MM211 GND! 326 178 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=7242  $PIN_XY=508,7326,478,7242,448,7326 $DEVICE_ID=1001
MM212 BL<0> WL<7> 326 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=6693  $PIN_XY=508,6696,478,6693,448,6696 $DEVICE_ID=1001
MM213 GND! 179 188 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=6318  $PIN_XY=508,6402,478,6318,448,6402 $DEVICE_ID=1001
MM214 BL<0> WL<6> 179 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=5769  $PIN_XY=508,5772,478,5769,448,5772 $DEVICE_ID=1001
MM215 GND! 189 172 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=5394  $PIN_XY=508,5478,478,5394,448,5478 $DEVICE_ID=1001
MM216 BL<0> WL<5> 189 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=4845  $PIN_XY=508,4848,478,4845,448,4848 $DEVICE_ID=1001
MM217 GND! 173 66 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=4470  $PIN_XY=508,4554,478,4470,448,4554 $DEVICE_ID=1001
MM218 178 WL<7> BLB<0> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=7329  $PIN_XY=340,7326,310,7329,280,7326 $DEVICE_ID=1001
MM219 326 178 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=6780  $PIN_XY=340,6696,310,6780,280,6696 $DEVICE_ID=1001
MM220 188 WL<6> BLB<0> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=6405  $PIN_XY=340,6402,310,6405,280,6402 $DEVICE_ID=1001
MM221 179 188 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=5856  $PIN_XY=340,5772,310,5856,280,5772 $DEVICE_ID=1001
MM222 172 WL<5> BLB<0> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=5481  $PIN_XY=340,5478,310,5481,280,5478 $DEVICE_ID=1001
MM223 189 172 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=4932  $PIN_XY=340,4848,310,4932,280,4848 $DEVICE_ID=1001
MM224 66 WL<4> BLB<0> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=4557  $PIN_XY=340,4554,310,4557,280,4554 $DEVICE_ID=1001
MM225 BL<15> WL<4> 249 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=3921  $PIN_XY=9076,3924,9046,3921,9016,3924 $DEVICE_ID=1001
MM226 GND! 159 148 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=3546  $PIN_XY=9076,3630,9046,3546,9016,3630 $DEVICE_ID=1001
MM227 BL<15> WL<3> 159 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=2997  $PIN_XY=9076,3000,9046,2997,9016,3000 $DEVICE_ID=1001
MM228 GND! 149 150 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=2622  $PIN_XY=9076,2706,9046,2622,9016,2706 $DEVICE_ID=1001
MM229 BL<15> WL<2> 149 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=2073  $PIN_XY=9076,2076,9046,2073,9016,2076 $DEVICE_ID=1001
MM230 GND! 151 168 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=1698  $PIN_XY=9076,1782,9046,1698,9016,1782 $DEVICE_ID=1001
MM231 BL<15> WL<1> 151 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=1149  $PIN_XY=9076,1152,9046,1149,9016,1152 $DEVICE_ID=1001
MM232 249 158 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=4008  $PIN_XY=8908,3924,8878,4008,8848,3924 $DEVICE_ID=1001
MM233 148 WL<3> BLB<15> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=3633  $PIN_XY=8908,3630,8878,3633,8848,3630 $DEVICE_ID=1001
MM234 159 148 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=3084  $PIN_XY=8908,3000,8878,3084,8848,3000 $DEVICE_ID=1001
MM235 150 WL<2> BLB<15> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=2709  $PIN_XY=8908,2706,8878,2709,8848,2706 $DEVICE_ID=1001
MM236 149 150 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=2160  $PIN_XY=8908,2076,8878,2160,8848,2076 $DEVICE_ID=1001
MM237 168 WL<1> BLB<15> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=1785  $PIN_XY=8908,1782,8878,1785,8848,1782 $DEVICE_ID=1001
MM238 151 168 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=1236  $PIN_XY=8908,1152,8878,1236,8848,1152 $DEVICE_ID=1001
MM239 BL<14> WL<4> 251 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=3921  $PIN_XY=8572,3924,8542,3921,8512,3924 $DEVICE_ID=1001
MM240 GND! 157 152 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=3546  $PIN_XY=8572,3630,8542,3546,8512,3630 $DEVICE_ID=1001
MM241 BL<14> WL<3> 157 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=2997  $PIN_XY=8572,3000,8542,2997,8512,3000 $DEVICE_ID=1001
MM242 GND! 153 154 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=2622  $PIN_XY=8572,2706,8542,2622,8512,2706 $DEVICE_ID=1001
MM243 BL<14> WL<2> 153 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=2073  $PIN_XY=8572,2076,8542,2073,8512,2076 $DEVICE_ID=1001
MM244 GND! 155 170 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=1698  $PIN_XY=8572,1782,8542,1698,8512,1782 $DEVICE_ID=1001
MM245 BL<14> WL<1> 155 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=1149  $PIN_XY=8572,1152,8542,1149,8512,1152 $DEVICE_ID=1001
MM246 251 156 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=4008  $PIN_XY=8404,3924,8374,4008,8344,3924 $DEVICE_ID=1001
MM247 152 WL<3> BLB<14> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=3633  $PIN_XY=8404,3630,8374,3633,8344,3630 $DEVICE_ID=1001
MM248 157 152 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=3084  $PIN_XY=8404,3000,8374,3084,8344,3000 $DEVICE_ID=1001
MM249 154 WL<2> BLB<14> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=2709  $PIN_XY=8404,2706,8374,2709,8344,2706 $DEVICE_ID=1001
MM250 153 154 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=2160  $PIN_XY=8404,2076,8374,2160,8344,2076 $DEVICE_ID=1001
MM251 170 WL<1> BLB<14> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=1785  $PIN_XY=8404,1782,8374,1785,8344,1782 $DEVICE_ID=1001
MM252 155 170 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=1236  $PIN_XY=8404,1152,8374,1236,8344,1152 $DEVICE_ID=1001
MM253 BL<13> WL<4> 247 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=3921  $PIN_XY=8068,3924,8038,3921,8008,3924 $DEVICE_ID=1001
MM254 GND! 161 144 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=3546  $PIN_XY=8068,3630,8038,3546,8008,3630 $DEVICE_ID=1001
MM255 BL<13> WL<3> 161 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=2997  $PIN_XY=8068,3000,8038,2997,8008,3000 $DEVICE_ID=1001
MM256 GND! 145 146 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=2622  $PIN_XY=8068,2706,8038,2622,8008,2706 $DEVICE_ID=1001
MM257 BL<13> WL<2> 145 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=2073  $PIN_XY=8068,2076,8038,2073,8008,2076 $DEVICE_ID=1001
MM258 GND! 147 166 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=1698  $PIN_XY=8068,1782,8038,1698,8008,1782 $DEVICE_ID=1001
MM259 BL<13> WL<1> 147 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=1149  $PIN_XY=8068,1152,8038,1149,8008,1152 $DEVICE_ID=1001
MM260 247 160 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=4008  $PIN_XY=7900,3924,7870,4008,7840,3924 $DEVICE_ID=1001
MM261 144 WL<3> BLB<13> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=3633  $PIN_XY=7900,3630,7870,3633,7840,3630 $DEVICE_ID=1001
MM262 161 144 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=3084  $PIN_XY=7900,3000,7870,3084,7840,3000 $DEVICE_ID=1001
MM263 146 WL<2> BLB<13> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=2709  $PIN_XY=7900,2706,7870,2709,7840,2706 $DEVICE_ID=1001
MM264 145 146 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=2160  $PIN_XY=7900,2076,7870,2160,7840,2076 $DEVICE_ID=1001
MM265 166 WL<1> BLB<13> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=1785  $PIN_XY=7900,1782,7870,1785,7840,1782 $DEVICE_ID=1001
MM266 147 166 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=1236  $PIN_XY=7900,1152,7870,1236,7840,1152 $DEVICE_ID=1001
MM267 BL<12> WL<4> 245 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=3921  $PIN_XY=7564,3924,7534,3921,7504,3924 $DEVICE_ID=1001
MM268 GND! 163 140 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=3546  $PIN_XY=7564,3630,7534,3546,7504,3630 $DEVICE_ID=1001
MM269 BL<12> WL<3> 163 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=2997  $PIN_XY=7564,3000,7534,2997,7504,3000 $DEVICE_ID=1001
MM270 GND! 141 142 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=2622  $PIN_XY=7564,2706,7534,2622,7504,2706 $DEVICE_ID=1001
MM271 BL<12> WL<2> 141 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=2073  $PIN_XY=7564,2076,7534,2073,7504,2076 $DEVICE_ID=1001
MM272 GND! 143 164 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=1698  $PIN_XY=7564,1782,7534,1698,7504,1782 $DEVICE_ID=1001
MM273 BL<12> WL<1> 143 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=1149  $PIN_XY=7564,1152,7534,1149,7504,1152 $DEVICE_ID=1001
MM274 245 162 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=4008  $PIN_XY=7396,3924,7366,4008,7336,3924 $DEVICE_ID=1001
MM275 140 WL<3> BLB<12> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=3633  $PIN_XY=7396,3630,7366,3633,7336,3630 $DEVICE_ID=1001
MM276 163 140 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=3084  $PIN_XY=7396,3000,7366,3084,7336,3000 $DEVICE_ID=1001
MM277 142 WL<2> BLB<12> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=2709  $PIN_XY=7396,2706,7366,2709,7336,2706 $DEVICE_ID=1001
MM278 141 142 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=2160  $PIN_XY=7396,2076,7366,2160,7336,2076 $DEVICE_ID=1001
MM279 164 WL<1> BLB<12> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=1785  $PIN_XY=7396,1782,7366,1785,7336,1782 $DEVICE_ID=1001
MM280 143 164 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=1236  $PIN_XY=7396,1152,7366,1236,7336,1152 $DEVICE_ID=1001
MM281 BL<11> WL<4> 229 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=3921  $PIN_XY=6724,3924,6694,3921,6664,3924 $DEVICE_ID=1001
MM282 GND! 131 120 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=3546  $PIN_XY=6724,3630,6694,3546,6664,3630 $DEVICE_ID=1001
MM283 BL<11> WL<3> 131 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=2997  $PIN_XY=6724,3000,6694,2997,6664,3000 $DEVICE_ID=1001
MM284 GND! 121 122 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=2622  $PIN_XY=6724,2706,6694,2622,6664,2706 $DEVICE_ID=1001
MM285 BL<11> WL<2> 121 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=2073  $PIN_XY=6724,2076,6694,2073,6664,2076 $DEVICE_ID=1001
MM286 GND! 123 136 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=1698  $PIN_XY=6724,1782,6694,1698,6664,1782 $DEVICE_ID=1001
MM287 BL<11> WL<1> 123 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=1149  $PIN_XY=6724,1152,6694,1149,6664,1152 $DEVICE_ID=1001
MM288 229 130 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=4008  $PIN_XY=6556,3924,6526,4008,6496,3924 $DEVICE_ID=1001
MM289 120 WL<3> BLB<11> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=3633  $PIN_XY=6556,3630,6526,3633,6496,3630 $DEVICE_ID=1001
MM290 131 120 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=3084  $PIN_XY=6556,3000,6526,3084,6496,3000 $DEVICE_ID=1001
MM291 122 WL<2> BLB<11> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=2709  $PIN_XY=6556,2706,6526,2709,6496,2706 $DEVICE_ID=1001
MM292 121 122 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=2160  $PIN_XY=6556,2076,6526,2160,6496,2076 $DEVICE_ID=1001
MM293 136 WL<1> BLB<11> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=1785  $PIN_XY=6556,1782,6526,1785,6496,1782 $DEVICE_ID=1001
MM294 123 136 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=1236  $PIN_XY=6556,1152,6526,1236,6496,1152 $DEVICE_ID=1001
MM295 BL<10> WL<4> 227 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=3921  $PIN_XY=6220,3924,6190,3921,6160,3924 $DEVICE_ID=1001
MM296 GND! 133 116 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=3546  $PIN_XY=6220,3630,6190,3546,6160,3630 $DEVICE_ID=1001
MM297 BL<10> WL<3> 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=2997  $PIN_XY=6220,3000,6190,2997,6160,3000 $DEVICE_ID=1001
MM298 GND! 117 118 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=2622  $PIN_XY=6220,2706,6190,2622,6160,2706 $DEVICE_ID=1001
MM299 BL<10> WL<2> 117 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=2073  $PIN_XY=6220,2076,6190,2073,6160,2076 $DEVICE_ID=1001
MM300 GND! 119 134 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=1698  $PIN_XY=6220,1782,6190,1698,6160,1782 $DEVICE_ID=1001
MM301 BL<10> WL<1> 119 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=1149  $PIN_XY=6220,1152,6190,1149,6160,1152 $DEVICE_ID=1001
MM302 227 132 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=4008  $PIN_XY=6052,3924,6022,4008,5992,3924 $DEVICE_ID=1001
MM303 116 WL<3> BLB<10> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=3633  $PIN_XY=6052,3630,6022,3633,5992,3630 $DEVICE_ID=1001
MM304 133 116 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=3084  $PIN_XY=6052,3000,6022,3084,5992,3000 $DEVICE_ID=1001
MM305 118 WL<2> BLB<10> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=2709  $PIN_XY=6052,2706,6022,2709,5992,2706 $DEVICE_ID=1001
MM306 117 118 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=2160  $PIN_XY=6052,2076,6022,2160,5992,2076 $DEVICE_ID=1001
MM307 134 WL<1> BLB<10> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=1785  $PIN_XY=6052,1782,6022,1785,5992,1782 $DEVICE_ID=1001
MM308 119 134 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=1236  $PIN_XY=6052,1152,6022,1236,5992,1152 $DEVICE_ID=1001
MM309 BL<9> WL<4> 231 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=3921  $PIN_XY=5716,3924,5686,3921,5656,3924 $DEVICE_ID=1001
MM310 GND! 129 124 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=3546  $PIN_XY=5716,3630,5686,3546,5656,3630 $DEVICE_ID=1001
MM311 BL<9> WL<3> 129 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=2997  $PIN_XY=5716,3000,5686,2997,5656,3000 $DEVICE_ID=1001
MM312 GND! 125 126 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=2622  $PIN_XY=5716,2706,5686,2622,5656,2706 $DEVICE_ID=1001
MM313 BL<9> WL<2> 125 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=2073  $PIN_XY=5716,2076,5686,2073,5656,2076 $DEVICE_ID=1001
MM314 GND! 127 138 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=1698  $PIN_XY=5716,1782,5686,1698,5656,1782 $DEVICE_ID=1001
MM315 BL<9> WL<1> 127 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=1149  $PIN_XY=5716,1152,5686,1149,5656,1152 $DEVICE_ID=1001
MM316 231 128 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=4008  $PIN_XY=5548,3924,5518,4008,5488,3924 $DEVICE_ID=1001
MM317 124 WL<3> BLB<9> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=3633  $PIN_XY=5548,3630,5518,3633,5488,3630 $DEVICE_ID=1001
MM318 129 124 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=3084  $PIN_XY=5548,3000,5518,3084,5488,3000 $DEVICE_ID=1001
MM319 126 WL<2> BLB<9> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=2709  $PIN_XY=5548,2706,5518,2709,5488,2706 $DEVICE_ID=1001
MM320 125 126 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=2160  $PIN_XY=5548,2076,5518,2160,5488,2076 $DEVICE_ID=1001
MM321 138 WL<1> BLB<9> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=1785  $PIN_XY=5548,1782,5518,1785,5488,1782 $DEVICE_ID=1001
MM322 127 138 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=1236  $PIN_XY=5548,1152,5518,1236,5488,1152 $DEVICE_ID=1001
MM323 BL<8> WL<4> 213 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=3921  $PIN_XY=5212,3924,5182,3921,5152,3924 $DEVICE_ID=1001
MM324 GND! 105 100 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=3546  $PIN_XY=5212,3630,5182,3546,5152,3630 $DEVICE_ID=1001
MM325 BL<8> WL<3> 105 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=2997  $PIN_XY=5212,3000,5182,2997,5152,3000 $DEVICE_ID=1001
MM326 GND! 101 102 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=2622  $PIN_XY=5212,2706,5182,2622,5152,2706 $DEVICE_ID=1001
MM327 BL<8> WL<2> 101 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=2073  $PIN_XY=5212,2076,5182,2073,5152,2076 $DEVICE_ID=1001
MM328 GND! 103 114 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=1698  $PIN_XY=5212,1782,5182,1698,5152,1782 $DEVICE_ID=1001
MM329 BL<8> WL<1> 103 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=1149  $PIN_XY=5212,1152,5182,1149,5152,1152 $DEVICE_ID=1001
MM330 213 104 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=4008  $PIN_XY=5044,3924,5014,4008,4984,3924 $DEVICE_ID=1001
MM331 100 WL<3> BLB<8> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=3633  $PIN_XY=5044,3630,5014,3633,4984,3630 $DEVICE_ID=1001
MM332 105 100 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=3084  $PIN_XY=5044,3000,5014,3084,4984,3000 $DEVICE_ID=1001
MM333 102 WL<2> BLB<8> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=2709  $PIN_XY=5044,2706,5014,2709,4984,2706 $DEVICE_ID=1001
MM334 101 102 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=2160  $PIN_XY=5044,2076,5014,2160,4984,2076 $DEVICE_ID=1001
MM335 114 WL<1> BLB<8> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=1785  $PIN_XY=5044,1782,5014,1785,4984,1782 $DEVICE_ID=1001
MM336 103 114 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=1236  $PIN_XY=5044,1152,5014,1236,4984,1152 $DEVICE_ID=1001
MM337 BL<7> WL<4> 211 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=3921  $PIN_XY=4372,3924,4342,3921,4312,3924 $DEVICE_ID=1001
MM338 GND! 107 96 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=3546  $PIN_XY=4372,3630,4342,3546,4312,3630 $DEVICE_ID=1001
MM339 BL<7> WL<3> 107 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=2997  $PIN_XY=4372,3000,4342,2997,4312,3000 $DEVICE_ID=1001
MM340 GND! 97 98 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=2622  $PIN_XY=4372,2706,4342,2622,4312,2706 $DEVICE_ID=1001
MM341 BL<7> WL<2> 97 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=2073  $PIN_XY=4372,2076,4342,2073,4312,2076 $DEVICE_ID=1001
MM342 GND! 99 112 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=1698  $PIN_XY=4372,1782,4342,1698,4312,1782 $DEVICE_ID=1001
MM343 BL<7> WL<1> 99 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=1149  $PIN_XY=4372,1152,4342,1149,4312,1152 $DEVICE_ID=1001
MM344 211 106 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=4008  $PIN_XY=4204,3924,4174,4008,4144,3924 $DEVICE_ID=1001
MM345 96 WL<3> BLB<7> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=3633  $PIN_XY=4204,3630,4174,3633,4144,3630 $DEVICE_ID=1001
MM346 107 96 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=3084  $PIN_XY=4204,3000,4174,3084,4144,3000 $DEVICE_ID=1001
MM347 98 WL<2> BLB<7> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=2709  $PIN_XY=4204,2706,4174,2709,4144,2706 $DEVICE_ID=1001
MM348 97 98 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=2160  $PIN_XY=4204,2076,4174,2160,4144,2076 $DEVICE_ID=1001
MM349 112 WL<1> BLB<7> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=1785  $PIN_XY=4204,1782,4174,1785,4144,1782 $DEVICE_ID=1001
MM350 99 112 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=1236  $PIN_XY=4204,1152,4174,1236,4144,1152 $DEVICE_ID=1001
MM351 BL<6> WL<4> 209 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=3921  $PIN_XY=3868,3924,3838,3921,3808,3924 $DEVICE_ID=1001
MM352 GND! 109 92 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=3546  $PIN_XY=3868,3630,3838,3546,3808,3630 $DEVICE_ID=1001
MM353 BL<6> WL<3> 109 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=2997  $PIN_XY=3868,3000,3838,2997,3808,3000 $DEVICE_ID=1001
MM354 GND! 93 94 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=2622  $PIN_XY=3868,2706,3838,2622,3808,2706 $DEVICE_ID=1001
MM355 BL<6> WL<2> 93 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=2073  $PIN_XY=3868,2076,3838,2073,3808,2076 $DEVICE_ID=1001
MM356 GND! 95 110 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=1698  $PIN_XY=3868,1782,3838,1698,3808,1782 $DEVICE_ID=1001
MM357 BL<6> WL<1> 95 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=1149  $PIN_XY=3868,1152,3838,1149,3808,1152 $DEVICE_ID=1001
MM358 209 108 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=4008  $PIN_XY=3700,3924,3670,4008,3640,3924 $DEVICE_ID=1001
MM359 92 WL<3> BLB<6> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=3633  $PIN_XY=3700,3630,3670,3633,3640,3630 $DEVICE_ID=1001
MM360 109 92 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=3084  $PIN_XY=3700,3000,3670,3084,3640,3000 $DEVICE_ID=1001
MM361 94 WL<2> BLB<6> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=2709  $PIN_XY=3700,2706,3670,2709,3640,2706 $DEVICE_ID=1001
MM362 93 94 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=2160  $PIN_XY=3700,2076,3670,2160,3640,2076 $DEVICE_ID=1001
MM363 110 WL<1> BLB<6> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=1785  $PIN_XY=3700,1782,3670,1785,3640,1782 $DEVICE_ID=1001
MM364 95 110 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=1236  $PIN_XY=3700,1152,3670,1236,3640,1152 $DEVICE_ID=1001
MM365 BL<5> WL<4> 193 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=3921  $PIN_XY=3364,3924,3334,3921,3304,3924 $DEVICE_ID=1001
MM366 GND! 83 72 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=3546  $PIN_XY=3364,3630,3334,3546,3304,3630 $DEVICE_ID=1001
MM367 BL<5> WL<3> 83 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=2997  $PIN_XY=3364,3000,3334,2997,3304,3000 $DEVICE_ID=1001
MM368 GND! 73 74 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=2622  $PIN_XY=3364,2706,3334,2622,3304,2706 $DEVICE_ID=1001
MM369 BL<5> WL<2> 73 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=2073  $PIN_XY=3364,2076,3334,2073,3304,2076 $DEVICE_ID=1001
MM370 GND! 75 86 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=1698  $PIN_XY=3364,1782,3334,1698,3304,1782 $DEVICE_ID=1001
MM371 BL<5> WL<1> 75 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=1149  $PIN_XY=3364,1152,3334,1149,3304,1152 $DEVICE_ID=1001
MM372 193 82 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=4008  $PIN_XY=3196,3924,3166,4008,3136,3924 $DEVICE_ID=1001
MM373 72 WL<3> BLB<5> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=3633  $PIN_XY=3196,3630,3166,3633,3136,3630 $DEVICE_ID=1001
MM374 83 72 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=3084  $PIN_XY=3196,3000,3166,3084,3136,3000 $DEVICE_ID=1001
MM375 74 WL<2> BLB<5> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=2709  $PIN_XY=3196,2706,3166,2709,3136,2706 $DEVICE_ID=1001
MM376 73 74 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=2160  $PIN_XY=3196,2076,3166,2160,3136,2076 $DEVICE_ID=1001
MM377 86 WL<1> BLB<5> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=1785  $PIN_XY=3196,1782,3166,1785,3136,1782 $DEVICE_ID=1001
MM378 75 86 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=1236  $PIN_XY=3196,1152,3166,1236,3136,1152 $DEVICE_ID=1001
MM379 BL<4> WL<4> 195 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=3921  $PIN_XY=2860,3924,2830,3921,2800,3924 $DEVICE_ID=1001
MM380 GND! 81 76 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=3546  $PIN_XY=2860,3630,2830,3546,2800,3630 $DEVICE_ID=1001
MM381 BL<4> WL<3> 81 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=2997  $PIN_XY=2860,3000,2830,2997,2800,3000 $DEVICE_ID=1001
MM382 GND! 77 78 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=2622  $PIN_XY=2860,2706,2830,2622,2800,2706 $DEVICE_ID=1001
MM383 BL<4> WL<2> 77 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=2073  $PIN_XY=2860,2076,2830,2073,2800,2076 $DEVICE_ID=1001
MM384 GND! 79 88 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=1698  $PIN_XY=2860,1782,2830,1698,2800,1782 $DEVICE_ID=1001
MM385 BL<4> WL<1> 79 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=1149  $PIN_XY=2860,1152,2830,1149,2800,1152 $DEVICE_ID=1001
MM386 195 80 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=4008  $PIN_XY=2692,3924,2662,4008,2632,3924 $DEVICE_ID=1001
MM387 76 WL<3> BLB<4> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=3633  $PIN_XY=2692,3630,2662,3633,2632,3630 $DEVICE_ID=1001
MM388 81 76 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=3084  $PIN_XY=2692,3000,2662,3084,2632,3000 $DEVICE_ID=1001
MM389 78 WL<2> BLB<4> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=2709  $PIN_XY=2692,2706,2662,2709,2632,2706 $DEVICE_ID=1001
MM390 77 78 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=2160  $PIN_XY=2692,2076,2662,2160,2632,2076 $DEVICE_ID=1001
MM391 88 WL<1> BLB<4> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=1785  $PIN_XY=2692,1782,2662,1785,2632,1782 $DEVICE_ID=1001
MM392 79 88 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=1236  $PIN_XY=2692,1152,2662,1236,2632,1152 $DEVICE_ID=1001
MM393 BL<3> WL<4> 191 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=3921  $PIN_XY=2020,3924,1990,3921,1960,3924 $DEVICE_ID=1001
MM394 GND! 91 70 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=3546  $PIN_XY=2020,3630,1990,3546,1960,3630 $DEVICE_ID=1001
MM395 BL<3> WL<3> 91 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=2997  $PIN_XY=2020,3000,1990,2997,1960,3000 $DEVICE_ID=1001
MM396 GND! 71 68 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=2622  $PIN_XY=2020,2706,1990,2622,1960,2706 $DEVICE_ID=1001
MM397 BL<3> WL<2> 71 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=2073  $PIN_XY=2020,2076,1990,2073,1960,2076 $DEVICE_ID=1001
MM398 GND! 69 84 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=1698  $PIN_XY=2020,1782,1990,1698,1960,1782 $DEVICE_ID=1001
MM399 BL<3> WL<1> 69 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=1149  $PIN_XY=2020,1152,1990,1149,1960,1152 $DEVICE_ID=1001
MM400 191 90 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=4008  $PIN_XY=1852,3924,1822,4008,1792,3924 $DEVICE_ID=1001
MM401 70 WL<3> BLB<3> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=3633  $PIN_XY=1852,3630,1822,3633,1792,3630 $DEVICE_ID=1001
MM402 91 70 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=3084  $PIN_XY=1852,3000,1822,3084,1792,3000 $DEVICE_ID=1001
MM403 68 WL<2> BLB<3> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=2709  $PIN_XY=1852,2706,1822,2709,1792,2706 $DEVICE_ID=1001
MM404 71 68 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=2160  $PIN_XY=1852,2076,1822,2160,1792,2076 $DEVICE_ID=1001
MM405 84 WL<1> BLB<3> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=1785  $PIN_XY=1852,1782,1822,1785,1792,1782 $DEVICE_ID=1001
MM406 69 84 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=1236  $PIN_XY=1852,1152,1822,1236,1792,1152 $DEVICE_ID=1001
MM407 BL<2> WL<4> 177 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=3921  $PIN_XY=1516,3924,1486,3921,1456,3924 $DEVICE_ID=1001
MM408 GND! 63 54 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=3546  $PIN_XY=1516,3630,1486,3546,1456,3630 $DEVICE_ID=1001
MM409 BL<2> WL<3> 63 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=2997  $PIN_XY=1516,3000,1486,2997,1456,3000 $DEVICE_ID=1001
MM410 GND! 55 52 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=2622  $PIN_XY=1516,2706,1486,2622,1456,2706 $DEVICE_ID=1001
MM411 BL<2> WL<2> 55 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=2073  $PIN_XY=1516,2076,1486,2073,1456,2076 $DEVICE_ID=1001
MM412 GND! 53 60 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=1698  $PIN_XY=1516,1782,1486,1698,1456,1782 $DEVICE_ID=1001
MM413 BL<2> WL<1> 53 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=1149  $PIN_XY=1516,1152,1486,1149,1456,1152 $DEVICE_ID=1001
MM414 177 62 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=4008  $PIN_XY=1348,3924,1318,4008,1288,3924 $DEVICE_ID=1001
MM415 54 WL<3> BLB<2> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=3633  $PIN_XY=1348,3630,1318,3633,1288,3630 $DEVICE_ID=1001
MM416 63 54 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=3084  $PIN_XY=1348,3000,1318,3084,1288,3000 $DEVICE_ID=1001
MM417 52 WL<2> BLB<2> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=2709  $PIN_XY=1348,2706,1318,2709,1288,2706 $DEVICE_ID=1001
MM418 55 52 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=2160  $PIN_XY=1348,2076,1318,2160,1288,2076 $DEVICE_ID=1001
MM419 60 WL<1> BLB<2> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=1785  $PIN_XY=1348,1782,1318,1785,1288,1782 $DEVICE_ID=1001
MM420 53 60 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=1236  $PIN_XY=1348,1152,1318,1236,1288,1152 $DEVICE_ID=1001
MM421 BL<1> WL<4> 175 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=3921  $PIN_XY=1012,3924,982,3921,952,3924 $DEVICE_ID=1001
MM422 GND! 65 50 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=3546  $PIN_XY=1012,3630,982,3546,952,3630 $DEVICE_ID=1001
MM423 BL<1> WL<3> 65 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=2997  $PIN_XY=1012,3000,982,2997,952,3000 $DEVICE_ID=1001
MM424 GND! 51 48 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=2622  $PIN_XY=1012,2706,982,2622,952,2706 $DEVICE_ID=1001
MM425 BL<1> WL<2> 51 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=2073  $PIN_XY=1012,2076,982,2073,952,2076 $DEVICE_ID=1001
MM426 GND! 49 58 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=1698  $PIN_XY=1012,1782,982,1698,952,1782 $DEVICE_ID=1001
MM427 BL<1> WL<1> 49 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=1149  $PIN_XY=1012,1152,982,1149,952,1152 $DEVICE_ID=1001
MM428 175 64 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=4008  $PIN_XY=844,3924,814,4008,784,3924 $DEVICE_ID=1001
MM429 50 WL<3> BLB<1> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=3633  $PIN_XY=844,3630,814,3633,784,3630 $DEVICE_ID=1001
MM430 65 50 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=3084  $PIN_XY=844,3000,814,3084,784,3000 $DEVICE_ID=1001
MM431 48 WL<2> BLB<1> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=2709  $PIN_XY=844,2706,814,2709,784,2706 $DEVICE_ID=1001
MM432 51 48 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=2160  $PIN_XY=844,2076,814,2160,784,2076 $DEVICE_ID=1001
MM433 58 WL<1> BLB<1> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=1785  $PIN_XY=844,1782,814,1785,784,1782 $DEVICE_ID=1001
MM434 49 58 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=1236  $PIN_XY=844,1152,814,1236,784,1152 $DEVICE_ID=1001
MM435 BL<0> WL<4> 173 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=3921  $PIN_XY=508,3924,478,3921,448,3924 $DEVICE_ID=1001
MM436 GND! 67 46 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=3546  $PIN_XY=508,3630,478,3546,448,3630 $DEVICE_ID=1001
MM437 BL<0> WL<3> 67 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=2997  $PIN_XY=508,3000,478,2997,448,3000 $DEVICE_ID=1001
MM438 GND! 47 44 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=2622  $PIN_XY=508,2706,478,2622,448,2706 $DEVICE_ID=1001
MM439 BL<0> WL<2> 47 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=2073  $PIN_XY=508,2076,478,2073,448,2076 $DEVICE_ID=1001
MM440 GND! 45 56 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=1698  $PIN_XY=508,1782,478,1698,448,1782 $DEVICE_ID=1001
MM441 BL<0> WL<1> 45 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=1149  $PIN_XY=508,1152,478,1149,448,1152 $DEVICE_ID=1001
MM442 173 66 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=4008  $PIN_XY=340,3924,310,4008,280,3924 $DEVICE_ID=1001
MM443 46 WL<3> BLB<0> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=3633  $PIN_XY=340,3630,310,3633,280,3630 $DEVICE_ID=1001
MM444 67 46 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=3084  $PIN_XY=340,3000,310,3084,280,3000 $DEVICE_ID=1001
MM445 44 WL<2> BLB<0> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=2709  $PIN_XY=340,2706,310,2709,280,2706 $DEVICE_ID=1001
MM446 47 44 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=2160  $PIN_XY=340,2076,310,2160,280,2076 $DEVICE_ID=1001
MM447 56 WL<1> BLB<0> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=1785  $PIN_XY=340,1782,310,1785,280,1782 $DEVICE_ID=1001
MM448 45 56 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=1236  $PIN_XY=340,1152,310,1236,280,1152 $DEVICE_ID=1001
MM449 GND! 169 317 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=774  $PIN_XY=9076,858,9046,774,9016,858 $DEVICE_ID=1001
MM450 BL<15> WL<0> 169 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=9046 $Y=225  $PIN_XY=9076,228,9046,225,9016,228 $DEVICE_ID=1001
MM451 317 WL<0> BLB<15> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=861  $PIN_XY=8908,858,8878,861,8848,858 $DEVICE_ID=1001
MM452 169 317 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8878 $Y=312  $PIN_XY=8908,228,8878,312,8848,228 $DEVICE_ID=1001
MM453 GND! 171 314 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=774  $PIN_XY=8572,858,8542,774,8512,858 $DEVICE_ID=1001
MM454 BL<14> WL<0> 171 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8542 $Y=225  $PIN_XY=8572,228,8542,225,8512,228 $DEVICE_ID=1001
MM455 314 WL<0> BLB<14> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=861  $PIN_XY=8404,858,8374,861,8344,858 $DEVICE_ID=1001
MM456 171 314 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=8374 $Y=312  $PIN_XY=8404,228,8374,312,8344,228 $DEVICE_ID=1001
MM457 GND! 167 320 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=774  $PIN_XY=8068,858,8038,774,8008,858 $DEVICE_ID=1001
MM458 BL<13> WL<0> 167 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=8038 $Y=225  $PIN_XY=8068,228,8038,225,8008,228 $DEVICE_ID=1001
MM459 320 WL<0> BLB<13> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=861  $PIN_XY=7900,858,7870,861,7840,858 $DEVICE_ID=1001
MM460 167 320 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7870 $Y=312  $PIN_XY=7900,228,7870,312,7840,228 $DEVICE_ID=1001
MM461 GND! 165 323 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=774  $PIN_XY=7564,858,7534,774,7504,858 $DEVICE_ID=1001
MM462 BL<12> WL<0> 165 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=7534 $Y=225  $PIN_XY=7564,228,7534,225,7504,228 $DEVICE_ID=1001
MM463 323 WL<0> BLB<12> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=861  $PIN_XY=7396,858,7366,861,7336,858 $DEVICE_ID=1001
MM464 165 323 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=7366 $Y=312  $PIN_XY=7396,228,7366,312,7336,228 $DEVICE_ID=1001
MM465 GND! 137 308 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=774  $PIN_XY=6724,858,6694,774,6664,858 $DEVICE_ID=1001
MM466 BL<11> WL<0> 137 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6694 $Y=225  $PIN_XY=6724,228,6694,225,6664,228 $DEVICE_ID=1001
MM467 308 WL<0> BLB<11> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=861  $PIN_XY=6556,858,6526,861,6496,858 $DEVICE_ID=1001
MM468 137 308 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6526 $Y=312  $PIN_XY=6556,228,6526,312,6496,228 $DEVICE_ID=1001
MM469 GND! 135 311 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=774  $PIN_XY=6220,858,6190,774,6160,858 $DEVICE_ID=1001
MM470 BL<10> WL<0> 135 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=6190 $Y=225  $PIN_XY=6220,228,6190,225,6160,228 $DEVICE_ID=1001
MM471 311 WL<0> BLB<10> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=861  $PIN_XY=6052,858,6022,861,5992,858 $DEVICE_ID=1001
MM472 135 311 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=6022 $Y=312  $PIN_XY=6052,228,6022,312,5992,228 $DEVICE_ID=1001
MM473 GND! 139 305 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=774  $PIN_XY=5716,858,5686,774,5656,858 $DEVICE_ID=1001
MM474 BL<9> WL<0> 139 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5686 $Y=225  $PIN_XY=5716,228,5686,225,5656,228 $DEVICE_ID=1001
MM475 305 WL<0> BLB<9> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=861  $PIN_XY=5548,858,5518,861,5488,858 $DEVICE_ID=1001
MM476 139 305 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5518 $Y=312  $PIN_XY=5548,228,5518,312,5488,228 $DEVICE_ID=1001
MM477 GND! 115 296 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=774  $PIN_XY=5212,858,5182,774,5152,858 $DEVICE_ID=1001
MM478 BL<8> WL<0> 115 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=5182 $Y=225  $PIN_XY=5212,228,5182,225,5152,228 $DEVICE_ID=1001
MM479 296 WL<0> BLB<8> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=861  $PIN_XY=5044,858,5014,861,4984,858 $DEVICE_ID=1001
MM480 115 296 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=5014 $Y=312  $PIN_XY=5044,228,5014,312,4984,228 $DEVICE_ID=1001
MM481 GND! 113 299 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=774  $PIN_XY=4372,858,4342,774,4312,858 $DEVICE_ID=1001
MM482 BL<7> WL<0> 113 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=4342 $Y=225  $PIN_XY=4372,228,4342,225,4312,228 $DEVICE_ID=1001
MM483 299 WL<0> BLB<7> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=861  $PIN_XY=4204,858,4174,861,4144,858 $DEVICE_ID=1001
MM484 113 299 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=4174 $Y=312  $PIN_XY=4204,228,4174,312,4144,228 $DEVICE_ID=1001
MM485 GND! 111 302 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=774  $PIN_XY=3868,858,3838,774,3808,858 $DEVICE_ID=1001
MM486 BL<6> WL<0> 111 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3838 $Y=225  $PIN_XY=3868,228,3838,225,3808,228 $DEVICE_ID=1001
MM487 302 WL<0> BLB<6> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=861  $PIN_XY=3700,858,3670,861,3640,858 $DEVICE_ID=1001
MM488 111 302 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3670 $Y=312  $PIN_XY=3700,228,3670,312,3640,228 $DEVICE_ID=1001
MM489 GND! 87 290 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=774  $PIN_XY=3364,858,3334,774,3304,858 $DEVICE_ID=1001
MM490 BL<5> WL<0> 87 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=3334 $Y=225  $PIN_XY=3364,228,3334,225,3304,228 $DEVICE_ID=1001
MM491 290 WL<0> BLB<5> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=861  $PIN_XY=3196,858,3166,861,3136,858 $DEVICE_ID=1001
MM492 87 290 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=3166 $Y=312  $PIN_XY=3196,228,3166,312,3136,228 $DEVICE_ID=1001
MM493 GND! 89 287 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=774  $PIN_XY=2860,858,2830,774,2800,858 $DEVICE_ID=1001
MM494 BL<4> WL<0> 89 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2830 $Y=225  $PIN_XY=2860,228,2830,225,2800,228 $DEVICE_ID=1001
MM495 287 WL<0> BLB<4> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=861  $PIN_XY=2692,858,2662,861,2632,858 $DEVICE_ID=1001
MM496 89 287 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2662 $Y=312  $PIN_XY=2692,228,2662,312,2632,228 $DEVICE_ID=1001
MM497 GND! 85 293 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=774  $PIN_XY=2020,858,1990,774,1960,858 $DEVICE_ID=1001
MM498 BL<3> WL<0> 85 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1990 $Y=225  $PIN_XY=2020,228,1990,225,1960,228 $DEVICE_ID=1001
MM499 293 WL<0> BLB<3> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=861  $PIN_XY=1852,858,1822,861,1792,858 $DEVICE_ID=1001
MM500 85 293 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1822 $Y=312  $PIN_XY=1852,228,1822,312,1792,228 $DEVICE_ID=1001
MM501 GND! 61 278 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=774  $PIN_XY=1516,858,1486,774,1456,858 $DEVICE_ID=1001
MM502 BL<2> WL<0> 61 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1486 $Y=225  $PIN_XY=1516,228,1486,225,1456,228 $DEVICE_ID=1001
MM503 278 WL<0> BLB<2> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=861  $PIN_XY=1348,858,1318,861,1288,858 $DEVICE_ID=1001
MM504 61 278 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1318 $Y=312  $PIN_XY=1348,228,1318,312,1288,228 $DEVICE_ID=1001
MM505 GND! 59 281 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=774  $PIN_XY=1012,858,982,774,952,858 $DEVICE_ID=1001
MM506 BL<1> WL<0> 59 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=982 $Y=225  $PIN_XY=1012,228,982,225,952,228 $DEVICE_ID=1001
MM507 281 WL<0> BLB<1> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=861  $PIN_XY=844,858,814,861,784,858 $DEVICE_ID=1001
MM508 59 281 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=814 $Y=312  $PIN_XY=844,228,814,312,784,228 $DEVICE_ID=1001
MM509 GND! 57 284 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=774  $PIN_XY=508,858,478,774,448,858 $DEVICE_ID=1001
MM510 BL<0> WL<0> 57 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=478 $Y=225  $PIN_XY=508,228,478,225,448,228 $DEVICE_ID=1001
MM511 284 WL<0> BLB<0> nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=861  $PIN_XY=340,858,310,861,280,858 $DEVICE_ID=1001
MM512 57 284 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=310 $Y=312  $PIN_XY=340,228,310,312,280,228 $DEVICE_ID=1001
XX246034E01 GND! VDD! 268 275 sram_filler $T=6804 7536 1 0 $X=6808 $Y=6946
XX246034E02 GND! VDD! 268 275 sram_filler $T=6804 6486 0 0 $X=6808 $Y=6486
XX246034E03 GND! VDD! 268 274 sram_filler $T=6804 4638 0 0 $X=6808 $Y=4638
XX246034E04 GND! VDD! 268 274 sram_filler $T=6804 5688 1 0 $X=6808 $Y=5098
XX246034E05 GND! VDD! 268 273 sram_filler $T=6804 4764 1 0 $X=6808 $Y=4174
XX246034E06 GND! VDD! 268 273 sram_filler $T=6804 3714 0 0 $X=6808 $Y=3714
XX246034E07 GND! VDD! 268 270 sram_filler $T=6804 18 0 0 $X=6808 $Y=18
XX246034E08 GND! VDD! 268 270 sram_filler $T=6804 1068 1 0 $X=6808 $Y=478
XX246034E09 GND! VDD! 268 269 sram_filler $T=6804 1992 1 0 $X=6808 $Y=1402
XX246034E010 GND! VDD! 268 269 sram_filler $T=6804 942 0 0 $X=6808 $Y=942
XX246034E011 GND! VDD! 268 272 sram_filler $T=6804 2790 0 0 $X=6808 $Y=2790
XX246034E012 GND! VDD! 268 272 sram_filler $T=6804 3840 1 0 $X=6808 $Y=3250
XX246034E013 GND! VDD! 268 271 sram_filler $T=6804 2916 1 0 $X=6808 $Y=2326
XX246034E014 GND! VDD! 268 271 sram_filler $T=6804 1866 0 0 $X=6808 $Y=1866
XX246034E015 GND! VDD! 268 276 sram_filler $T=6804 5562 0 0 $X=6808 $Y=5562
XX246034E016 GND! VDD! 268 276 sram_filler $T=6804 6612 1 0 $X=6808 $Y=6022
XX246034E017 GND! VDD! 268 270 sram_filler $T=4452 18 0 0 $X=4455 $Y=18
XX246034E018 GND! VDD! 268 270 sram_filler $T=4452 1068 1 0 $X=4455 $Y=478
XX246034E019 GND! VDD! 268 273 sram_filler $T=4452 3714 0 0 $X=4455 $Y=3714
XX246034E020 GND! VDD! 268 273 sram_filler $T=4452 4764 1 0 $X=4455 $Y=4174
XX246034E021 GND! VDD! 268 274 sram_filler $T=4452 5688 1 0 $X=4455 $Y=5098
XX246034E022 GND! VDD! 268 274 sram_filler $T=4452 4638 0 0 $X=4455 $Y=4638
XX246034E023 GND! VDD! 268 275 sram_filler $T=4452 6486 0 0 $X=4455 $Y=6486
XX246034E024 GND! VDD! 268 275 sram_filler $T=4452 7536 1 0 $X=4455 $Y=6946
XX246034E025 GND! VDD! 268 276 sram_filler $T=4452 6612 1 0 $X=4455 $Y=6022
XX246034E026 GND! VDD! 268 276 sram_filler $T=4452 5562 0 0 $X=4455 $Y=5562
XX246034E027 GND! VDD! 268 271 sram_filler $T=4452 1866 0 0 $X=4455 $Y=1866
XX246034E028 GND! VDD! 268 271 sram_filler $T=4452 2916 1 0 $X=4455 $Y=2326
XX246034E029 GND! VDD! 268 272 sram_filler $T=4452 3840 1 0 $X=4455 $Y=3250
XX246034E030 GND! VDD! 268 272 sram_filler $T=4452 2790 0 0 $X=4455 $Y=2790
XX246034E031 GND! VDD! 268 269 sram_filler $T=4452 942 0 0 $X=4455 $Y=942
XX246034E032 GND! VDD! 268 269 sram_filler $T=4452 1992 1 0 $X=4455 $Y=1402
XX246034E033 GND! VDD! 268 273 sram_filler $T=2100 3714 0 0 $X=2104 $Y=3714
XX246034E034 GND! VDD! 268 273 sram_filler $T=2100 4764 1 0 $X=2104 $Y=4174
XX246034E035 GND! VDD! 268 274 sram_filler $T=2100 5688 1 0 $X=2104 $Y=5098
XX246034E036 GND! VDD! 268 274 sram_filler $T=2100 4638 0 0 $X=2104 $Y=4638
XX246034E037 GND! VDD! 268 275 sram_filler $T=2100 6486 0 0 $X=2104 $Y=6486
XX246034E038 GND! VDD! 268 275 sram_filler $T=2100 7536 1 0 $X=2104 $Y=6946
XX246034E039 GND! VDD! 268 276 sram_filler $T=2100 6612 1 0 $X=2104 $Y=6022
XX246034E040 GND! VDD! 268 276 sram_filler $T=2100 5562 0 0 $X=2104 $Y=5562
XX246034E041 GND! VDD! 268 271 sram_filler $T=2100 1866 0 0 $X=2104 $Y=1866
XX246034E042 GND! VDD! 268 271 sram_filler $T=2100 2916 1 0 $X=2104 $Y=2326
XX246034E043 GND! VDD! 268 272 sram_filler $T=2100 3840 1 0 $X=2104 $Y=3250
XX246034E044 GND! VDD! 268 272 sram_filler $T=2100 2790 0 0 $X=2104 $Y=2790
XX246034E045 GND! VDD! 268 269 sram_filler $T=2100 942 0 0 $X=2104 $Y=942
XX246034E046 GND! VDD! 268 269 sram_filler $T=2100 1992 1 0 $X=2104 $Y=1402
XX246034E047 GND! VDD! 268 270 sram_filler $T=2100 1068 1 0 $X=2104 $Y=478
XX246034E048 GND! VDD! 268 270 sram_filler $T=2100 18 0 0 $X=2104 $Y=18
XX246034E049 GND! VDD! GND! BLB<0> 173 66 BL<0> WL<4> WL<3> 172 67 
+	WL<5> 268 268 273 sram_6t $T=112 3714 0 0 $X=88 $Y=3714
XX246034E050 GND! VDD! GND! BLB<1> 175 64 BL<1> WL<4> WL<3> 174 65 
+	WL<5> 268 268 273 sram_6t $T=616 3714 0 0 $X=592 $Y=3714
XX246034E051 GND! VDD! GND! BLB<3> 191 90 BL<3> WL<4> WL<3> 190 91 
+	WL<5> 268 268 273 sram_6t $T=1624 3714 0 0 $X=1600 $Y=3714
XX246034E052 GND! VDD! GND! BLB<2> 177 62 BL<2> WL<4> WL<3> 176 63 
+	WL<5> 268 268 273 sram_6t $T=1120 3714 0 0 $X=1096 $Y=3714
XX246034E053 GND! VDD! GND! BLB<6> 209 108 BL<6> WL<4> WL<3> 208 109 
+	WL<5> 268 268 273 sram_6t $T=3472 3714 0 0 $X=3448 $Y=3714
XX246034E054 GND! VDD! GND! BLB<7> 211 106 BL<7> WL<4> WL<3> 210 107 
+	WL<5> 268 268 273 sram_6t $T=3976 3714 0 0 $X=3952 $Y=3714
XX246034E055 GND! VDD! GND! BLB<5> 193 82 BL<5> WL<4> WL<3> 192 83 
+	WL<5> 268 268 273 sram_6t $T=2968 3714 0 0 $X=2944 $Y=3714
XX246034E056 GND! VDD! GND! BLB<4> 195 80 BL<4> WL<4> WL<3> 194 81 
+	WL<5> 268 268 273 sram_6t $T=2464 3714 0 0 $X=2440 $Y=3714
XX246034E057 GND! VDD! GND! BLB<12> 245 162 BL<12> WL<4> WL<3> 244 163 
+	WL<5> 268 268 273 sram_6t $T=7168 3714 0 0 $X=7144 $Y=3714
XX246034E058 GND! VDD! GND! BLB<13> 247 160 BL<13> WL<4> WL<3> 246 161 
+	WL<5> 268 268 273 sram_6t $T=7672 3714 0 0 $X=7648 $Y=3714
XX246034E059 GND! VDD! GND! BLB<15> 249 158 BL<15> WL<4> WL<3> 248 159 
+	WL<5> 268 268 273 sram_6t $T=8680 3714 0 0 $X=8656 $Y=3714
XX246034E060 GND! VDD! GND! BLB<14> 251 156 BL<14> WL<4> WL<3> 250 157 
+	WL<5> 268 268 273 sram_6t $T=8176 3714 0 0 $X=8152 $Y=3714
XX246034E061 GND! VDD! GND! BLB<0> 326 178 BL<0> WL<7> WL<6> 325 179 
+	327 268 268 275 sram_6t $T=112 6486 0 0 $X=88 $Y=6486
XX246034E062 GND! VDD! GND! BLB<1> 329 180 BL<1> WL<7> WL<6> 328 181 
+	330 268 268 275 sram_6t $T=616 6486 0 0 $X=592 $Y=6486
XX246034E063 GND! VDD! GND! BLB<10> 227 132 BL<10> WL<4> WL<3> 226 133 
+	WL<5> 268 268 273 sram_6t $T=5824 3714 0 0 $X=5800 $Y=3714
XX246034E064 GND! VDD! GND! BLB<11> 229 130 BL<11> WL<4> WL<3> 228 131 
+	WL<5> 268 268 273 sram_6t $T=6328 3714 0 0 $X=6304 $Y=3714
XX246034E065 GND! VDD! GND! BLB<9> 231 128 BL<9> WL<4> WL<3> 230 129 
+	WL<5> 268 268 273 sram_6t $T=5320 3714 0 0 $X=5296 $Y=3714
XX246034E066 GND! VDD! GND! BLB<8> 213 104 BL<8> WL<4> WL<3> 212 105 
+	WL<5> 268 268 273 sram_6t $T=4816 3714 0 0 $X=4792 $Y=3714
XX246034E067 GND! VDD! GND! BLB<8> 215 212 BL<8> WL<5> WL<4> 214 213 
+	WL<6> 268 268 274 sram_6t $T=4816 4638 0 0 $X=4792 $Y=4638
XX246034E068 GND! VDD! GND! BLB<9> 233 230 BL<9> WL<5> WL<4> 232 231 
+	WL<6> 268 268 274 sram_6t $T=5320 4638 0 0 $X=5296 $Y=4638
XX246034E069 GND! VDD! GND! BLB<11> 235 228 BL<11> WL<5> WL<4> 234 229 
+	WL<6> 268 268 274 sram_6t $T=6328 4638 0 0 $X=6304 $Y=4638
XX246034E070 GND! VDD! GND! BLB<10> 237 226 BL<10> WL<5> WL<4> 236 227 
+	WL<6> 268 268 274 sram_6t $T=5824 4638 0 0 $X=5800 $Y=4638
XX246034E071 GND! VDD! GND! BLB<2> 332 182 BL<2> WL<7> WL<6> 331 183 
+	333 268 268 275 sram_6t $T=1120 6486 0 0 $X=1096 $Y=6486
XX246034E072 GND! VDD! GND! BLB<3> 335 196 BL<3> WL<7> WL<6> 334 197 
+	336 268 268 275 sram_6t $T=1624 6486 0 0 $X=1600 $Y=6486
XX246034E073 GND! VDD! GND! BLB<14> 253 250 BL<14> WL<5> WL<4> 252 251 
+	WL<6> 268 268 274 sram_6t $T=8176 4638 0 0 $X=8152 $Y=4638
XX246034E074 GND! VDD! GND! BLB<15> 255 248 BL<15> WL<5> WL<4> 254 249 
+	WL<6> 268 268 274 sram_6t $T=8680 4638 0 0 $X=8656 $Y=4638
XX246034E075 GND! VDD! GND! BLB<13> 257 246 BL<13> WL<5> WL<4> 256 247 
+	WL<6> 268 268 274 sram_6t $T=7672 4638 0 0 $X=7648 $Y=4638
XX246034E076 GND! VDD! GND! BLB<12> 259 244 BL<12> WL<5> WL<4> 258 245 
+	WL<6> 268 268 274 sram_6t $T=7168 4638 0 0 $X=7144 $Y=4638
XX246034E077 GND! VDD! GND! BLB<4> 199 194 BL<4> WL<5> WL<4> 198 195 
+	WL<6> 268 268 274 sram_6t $T=2464 4638 0 0 $X=2440 $Y=4638
XX246034E078 GND! VDD! GND! BLB<5> 201 192 BL<5> WL<5> WL<4> 200 193 
+	WL<6> 268 268 274 sram_6t $T=2968 4638 0 0 $X=2944 $Y=4638
XX246034E079 GND! VDD! GND! BLB<7> 217 210 BL<7> WL<5> WL<4> 216 211 
+	WL<6> 268 268 274 sram_6t $T=3976 4638 0 0 $X=3952 $Y=4638
XX246034E080 GND! VDD! GND! BLB<6> 219 208 BL<6> WL<5> WL<4> 218 209 
+	WL<6> 268 268 274 sram_6t $T=3472 4638 0 0 $X=3448 $Y=4638
XX246034E081 GND! VDD! GND! BLB<2> 185 176 BL<2> WL<5> WL<4> 184 177 
+	WL<6> 268 268 274 sram_6t $T=1120 4638 0 0 $X=1096 $Y=4638
XX246034E082 GND! VDD! GND! BLB<3> 203 190 BL<3> WL<5> WL<4> 202 191 
+	WL<6> 268 268 274 sram_6t $T=1624 4638 0 0 $X=1600 $Y=4638
XX246034E083 GND! VDD! GND! BLB<1> 187 174 BL<1> WL<5> WL<4> 186 175 
+	WL<6> 268 268 274 sram_6t $T=616 4638 0 0 $X=592 $Y=4638
XX246034E084 GND! VDD! GND! BLB<0> 189 172 BL<0> WL<5> WL<4> 188 173 
+	WL<6> 268 268 274 sram_6t $T=112 4638 0 0 $X=88 $Y=4638
XX246034E085 GND! VDD! GND! BLB<6> 344 220 BL<6> WL<7> WL<6> 343 221 
+	345 268 268 275 sram_6t $T=3472 6486 0 0 $X=3448 $Y=6486
XX246034E086 GND! VDD! GND! BLB<7> 347 222 BL<7> WL<7> WL<6> 346 223 
+	348 268 268 275 sram_6t $T=3976 6486 0 0 $X=3952 $Y=6486
XX246034E087 GND! VDD! GND! BLB<5> 338 204 BL<5> WL<7> WL<6> 337 205 
+	339 268 268 275 sram_6t $T=2968 6486 0 0 $X=2944 $Y=6486
XX246034E088 GND! VDD! GND! BLB<4> 341 206 BL<4> WL<7> WL<6> 340 207 
+	342 268 268 275 sram_6t $T=2464 6486 0 0 $X=2440 $Y=6486
XX246034E089 GND! VDD! GND! BLB<12> 362 260 BL<12> WL<7> WL<6> 361 261 
+	363 268 268 275 sram_6t $T=7168 6486 0 0 $X=7144 $Y=6486
XX246034E090 GND! VDD! GND! BLB<13> 365 262 BL<13> WL<7> WL<6> 364 263 
+	366 268 268 275 sram_6t $T=7672 6486 0 0 $X=7648 $Y=6486
XX246034E091 GND! VDD! GND! BLB<15> 368 264 BL<15> WL<7> WL<6> 367 265 
+	369 268 268 275 sram_6t $T=8680 6486 0 0 $X=8656 $Y=6486
XX246034E092 GND! VDD! GND! BLB<14> 371 266 BL<14> WL<7> WL<6> 370 267 
+	372 268 268 275 sram_6t $T=8176 6486 0 0 $X=8152 $Y=6486
XX246034E093 GND! VDD! GND! BLB<10> 353 238 BL<10> WL<7> WL<6> 352 239 
+	354 268 268 275 sram_6t $T=5824 6486 0 0 $X=5800 $Y=6486
XX246034E094 GND! VDD! GND! BLB<11> 356 240 BL<11> WL<7> WL<6> 355 241 
+	357 268 268 275 sram_6t $T=6328 6486 0 0 $X=6304 $Y=6486
XX246034E095 GND! VDD! GND! BLB<9> 359 242 BL<9> WL<7> WL<6> 358 243 
+	360 268 268 275 sram_6t $T=5320 6486 0 0 $X=5296 $Y=6486
XX246034E096 GND! VDD! GND! BLB<8> 350 224 BL<8> WL<7> WL<6> 349 225 
+	351 268 268 275 sram_6t $T=4816 6486 0 0 $X=4792 $Y=6486
XX246034E097 GND! VDD! GND! BLB<8> 225 214 BL<8> WL<6> WL<5> 224 215 
+	WL<7> 268 268 276 sram_6t $T=4816 5562 0 0 $X=4792 $Y=5562
XX246034E098 GND! VDD! GND! BLB<9> 243 232 BL<9> WL<6> WL<5> 242 233 
+	WL<7> 268 268 276 sram_6t $T=5320 5562 0 0 $X=5296 $Y=5562
XX246034E099 GND! VDD! GND! BLB<11> 241 234 BL<11> WL<6> WL<5> 240 235 
+	WL<7> 268 268 276 sram_6t $T=6328 5562 0 0 $X=6304 $Y=5562
XX246034E0100 GND! VDD! GND! BLB<10> 239 236 BL<10> WL<6> WL<5> 238 237 
+	WL<7> 268 268 276 sram_6t $T=5824 5562 0 0 $X=5800 $Y=5562
XX246034E0101 GND! VDD! GND! BLB<14> 267 252 BL<14> WL<6> WL<5> 266 253 
+	WL<7> 268 268 276 sram_6t $T=8176 5562 0 0 $X=8152 $Y=5562
XX246034E0102 GND! VDD! GND! BLB<15> 265 254 BL<15> WL<6> WL<5> 264 255 
+	WL<7> 268 268 276 sram_6t $T=8680 5562 0 0 $X=8656 $Y=5562
XX246034E0103 GND! VDD! GND! BLB<13> 263 256 BL<13> WL<6> WL<5> 262 257 
+	WL<7> 268 268 276 sram_6t $T=7672 5562 0 0 $X=7648 $Y=5562
XX246034E0104 GND! VDD! GND! BLB<12> 261 258 BL<12> WL<6> WL<5> 260 259 
+	WL<7> 268 268 276 sram_6t $T=7168 5562 0 0 $X=7144 $Y=5562
XX246034E0105 GND! VDD! GND! BLB<4> 207 198 BL<4> WL<6> WL<5> 206 199 
+	WL<7> 268 268 276 sram_6t $T=2464 5562 0 0 $X=2440 $Y=5562
XX246034E0106 GND! VDD! GND! BLB<5> 205 200 BL<5> WL<6> WL<5> 204 201 
+	WL<7> 268 268 276 sram_6t $T=2968 5562 0 0 $X=2944 $Y=5562
XX246034E0107 GND! VDD! GND! BLB<7> 223 216 BL<7> WL<6> WL<5> 222 217 
+	WL<7> 268 268 276 sram_6t $T=3976 5562 0 0 $X=3952 $Y=5562
XX246034E0108 GND! VDD! GND! BLB<6> 221 218 BL<6> WL<6> WL<5> 220 219 
+	WL<7> 268 268 276 sram_6t $T=3472 5562 0 0 $X=3448 $Y=5562
XX246034E0109 GND! VDD! GND! BLB<2> 183 184 BL<2> WL<6> WL<5> 182 185 
+	WL<7> 268 268 276 sram_6t $T=1120 5562 0 0 $X=1096 $Y=5562
XX246034E0110 GND! VDD! GND! BLB<3> 197 202 BL<3> WL<6> WL<5> 196 203 
+	WL<7> 268 268 276 sram_6t $T=1624 5562 0 0 $X=1600 $Y=5562
XX246034E0111 GND! VDD! GND! BLB<1> 181 186 BL<1> WL<6> WL<5> 180 187 
+	WL<7> 268 268 276 sram_6t $T=616 5562 0 0 $X=592 $Y=5562
XX246034E0112 GND! VDD! GND! BLB<0> 179 188 BL<0> WL<6> WL<5> 178 189 
+	WL<7> 268 268 276 sram_6t $T=112 5562 0 0 $X=88 $Y=5562
XX246034E0113 GND! VDD! GND! BLB<0> 47 44 BL<0> WL<2> WL<1> 46 45 
+	WL<3> 268 268 271 sram_6t $T=112 1866 0 0 $X=88 $Y=1866
XX246034E0114 GND! VDD! GND! BLB<1> 51 48 BL<1> WL<2> WL<1> 50 49 
+	WL<3> 268 268 271 sram_6t $T=616 1866 0 0 $X=592 $Y=1866
XX246034E0115 GND! VDD! GND! BLB<3> 71 68 BL<3> WL<2> WL<1> 70 69 
+	WL<3> 268 268 271 sram_6t $T=1624 1866 0 0 $X=1600 $Y=1866
XX246034E0116 GND! VDD! GND! BLB<2> 55 52 BL<2> WL<2> WL<1> 54 53 
+	WL<3> 268 268 271 sram_6t $T=1120 1866 0 0 $X=1096 $Y=1866
XX246034E0117 GND! VDD! GND! BLB<6> 93 94 BL<6> WL<2> WL<1> 92 95 
+	WL<3> 268 268 271 sram_6t $T=3472 1866 0 0 $X=3448 $Y=1866
XX246034E0118 GND! VDD! GND! BLB<7> 97 98 BL<7> WL<2> WL<1> 96 99 
+	WL<3> 268 268 271 sram_6t $T=3976 1866 0 0 $X=3952 $Y=1866
XX246034E0119 GND! VDD! GND! BLB<5> 73 74 BL<5> WL<2> WL<1> 72 75 
+	WL<3> 268 268 271 sram_6t $T=2968 1866 0 0 $X=2944 $Y=1866
XX246034E0120 GND! VDD! GND! BLB<4> 77 78 BL<4> WL<2> WL<1> 76 79 
+	WL<3> 268 268 271 sram_6t $T=2464 1866 0 0 $X=2440 $Y=1866
XX246034E0121 GND! VDD! GND! BLB<12> 141 142 BL<12> WL<2> WL<1> 140 143 
+	WL<3> 268 268 271 sram_6t $T=7168 1866 0 0 $X=7144 $Y=1866
XX246034E0122 GND! VDD! GND! BLB<13> 145 146 BL<13> WL<2> WL<1> 144 147 
+	WL<3> 268 268 271 sram_6t $T=7672 1866 0 0 $X=7648 $Y=1866
XX246034E0123 GND! VDD! GND! BLB<15> 149 150 BL<15> WL<2> WL<1> 148 151 
+	WL<3> 268 268 271 sram_6t $T=8680 1866 0 0 $X=8656 $Y=1866
XX246034E0124 GND! VDD! GND! BLB<14> 153 154 BL<14> WL<2> WL<1> 152 155 
+	WL<3> 268 268 271 sram_6t $T=8176 1866 0 0 $X=8152 $Y=1866
XX246034E0125 GND! VDD! GND! BLB<10> 117 118 BL<10> WL<2> WL<1> 116 119 
+	WL<3> 268 268 271 sram_6t $T=5824 1866 0 0 $X=5800 $Y=1866
XX246034E0126 GND! VDD! GND! BLB<11> 121 122 BL<11> WL<2> WL<1> 120 123 
+	WL<3> 268 268 271 sram_6t $T=6328 1866 0 0 $X=6304 $Y=1866
XX246034E0127 GND! VDD! GND! BLB<9> 125 126 BL<9> WL<2> WL<1> 124 127 
+	WL<3> 268 268 271 sram_6t $T=5320 1866 0 0 $X=5296 $Y=1866
XX246034E0128 GND! VDD! GND! BLB<8> 101 102 BL<8> WL<2> WL<1> 100 103 
+	WL<3> 268 268 271 sram_6t $T=4816 1866 0 0 $X=4792 $Y=1866
XX246034E0129 GND! VDD! GND! BLB<8> 105 100 BL<8> WL<3> WL<2> 104 101 
+	WL<4> 268 268 272 sram_6t $T=4816 2790 0 0 $X=4792 $Y=2790
XX246034E0130 GND! VDD! GND! BLB<9> 129 124 BL<9> WL<3> WL<2> 128 125 
+	WL<4> 268 268 272 sram_6t $T=5320 2790 0 0 $X=5296 $Y=2790
XX246034E0131 GND! VDD! GND! BLB<11> 131 120 BL<11> WL<3> WL<2> 130 121 
+	WL<4> 268 268 272 sram_6t $T=6328 2790 0 0 $X=6304 $Y=2790
XX246034E0132 GND! VDD! GND! BLB<10> 133 116 BL<10> WL<3> WL<2> 132 117 
+	WL<4> 268 268 272 sram_6t $T=5824 2790 0 0 $X=5800 $Y=2790
XX246034E0133 GND! VDD! GND! BLB<14> 157 152 BL<14> WL<3> WL<2> 156 153 
+	WL<4> 268 268 272 sram_6t $T=8176 2790 0 0 $X=8152 $Y=2790
XX246034E0134 GND! VDD! GND! BLB<15> 159 148 BL<15> WL<3> WL<2> 158 149 
+	WL<4> 268 268 272 sram_6t $T=8680 2790 0 0 $X=8656 $Y=2790
XX246034E0135 GND! VDD! GND! BLB<13> 161 144 BL<13> WL<3> WL<2> 160 145 
+	WL<4> 268 268 272 sram_6t $T=7672 2790 0 0 $X=7648 $Y=2790
XX246034E0136 GND! VDD! GND! BLB<12> 163 140 BL<12> WL<3> WL<2> 162 141 
+	WL<4> 268 268 272 sram_6t $T=7168 2790 0 0 $X=7144 $Y=2790
XX246034E0137 GND! VDD! GND! BLB<4> 81 76 BL<4> WL<3> WL<2> 80 77 
+	WL<4> 268 268 272 sram_6t $T=2464 2790 0 0 $X=2440 $Y=2790
XX246034E0138 GND! VDD! GND! BLB<5> 83 72 BL<5> WL<3> WL<2> 82 73 
+	WL<4> 268 268 272 sram_6t $T=2968 2790 0 0 $X=2944 $Y=2790
XX246034E0139 GND! VDD! GND! BLB<7> 107 96 BL<7> WL<3> WL<2> 106 97 
+	WL<4> 268 268 272 sram_6t $T=3976 2790 0 0 $X=3952 $Y=2790
XX246034E0140 GND! VDD! GND! BLB<6> 109 92 BL<6> WL<3> WL<2> 108 93 
+	WL<4> 268 268 272 sram_6t $T=3472 2790 0 0 $X=3448 $Y=2790
XX246034E0141 GND! VDD! GND! BLB<0> 45 56 BL<0> WL<1> WL<0> 44 57 
+	WL<2> 268 268 269 sram_6t $T=112 942 0 0 $X=88 $Y=942
XX246034E0142 GND! VDD! GND! BLB<1> 49 58 BL<1> WL<1> WL<0> 48 59 
+	WL<2> 268 268 269 sram_6t $T=616 942 0 0 $X=592 $Y=942
XX246034E0143 GND! VDD! GND! BLB<3> 69 84 BL<3> WL<1> WL<0> 68 85 
+	WL<2> 268 268 269 sram_6t $T=1624 942 0 0 $X=1600 $Y=942
XX246034E0144 GND! VDD! GND! BLB<2> 53 60 BL<2> WL<1> WL<0> 52 61 
+	WL<2> 268 268 269 sram_6t $T=1120 942 0 0 $X=1096 $Y=942
XX246034E0145 GND! VDD! GND! BLB<6> 95 110 BL<6> WL<1> WL<0> 94 111 
+	WL<2> 268 268 269 sram_6t $T=3472 942 0 0 $X=3448 $Y=942
XX246034E0146 GND! VDD! GND! BLB<7> 99 112 BL<7> WL<1> WL<0> 98 113 
+	WL<2> 268 268 269 sram_6t $T=3976 942 0 0 $X=3952 $Y=942
XX246034E0147 GND! VDD! GND! BLB<5> 75 86 BL<5> WL<1> WL<0> 74 87 
+	WL<2> 268 268 269 sram_6t $T=2968 942 0 0 $X=2944 $Y=942
XX246034E0148 GND! VDD! GND! BLB<4> 79 88 BL<4> WL<1> WL<0> 78 89 
+	WL<2> 268 268 269 sram_6t $T=2464 942 0 0 $X=2440 $Y=942
XX246034E0149 GND! VDD! GND! BLB<12> 143 164 BL<12> WL<1> WL<0> 142 165 
+	WL<2> 268 268 269 sram_6t $T=7168 942 0 0 $X=7144 $Y=942
XX246034E0150 GND! VDD! GND! BLB<13> 147 166 BL<13> WL<1> WL<0> 146 167 
+	WL<2> 268 268 269 sram_6t $T=7672 942 0 0 $X=7648 $Y=942
XX246034E0151 GND! VDD! GND! BLB<15> 151 168 BL<15> WL<1> WL<0> 150 169 
+	WL<2> 268 268 269 sram_6t $T=8680 942 0 0 $X=8656 $Y=942
XX246034E0152 GND! VDD! GND! BLB<14> 155 170 BL<14> WL<1> WL<0> 154 171 
+	WL<2> 268 268 269 sram_6t $T=8176 942 0 0 $X=8152 $Y=942
XX246034E0153 GND! VDD! GND! BLB<3> 91 70 BL<3> WL<3> WL<2> 90 71 
+	WL<4> 268 268 272 sram_6t $T=1624 2790 0 0 $X=1600 $Y=2790
XX246034E0154 GND! VDD! GND! BLB<2> 63 54 BL<2> WL<3> WL<2> 62 55 
+	WL<4> 268 268 272 sram_6t $T=1120 2790 0 0 $X=1096 $Y=2790
XX246034E0155 GND! VDD! GND! BLB<10> 119 134 BL<10> WL<1> WL<0> 118 135 
+	WL<2> 268 268 269 sram_6t $T=5824 942 0 0 $X=5800 $Y=942
XX246034E0156 GND! VDD! GND! BLB<11> 123 136 BL<11> WL<1> WL<0> 122 137 
+	WL<2> 268 268 269 sram_6t $T=6328 942 0 0 $X=6304 $Y=942
XX246034E0157 GND! VDD! GND! BLB<9> 127 138 BL<9> WL<1> WL<0> 126 139 
+	WL<2> 268 268 269 sram_6t $T=5320 942 0 0 $X=5296 $Y=942
XX246034E0158 GND! VDD! GND! BLB<8> 103 114 BL<8> WL<1> WL<0> 102 115 
+	WL<2> 268 268 269 sram_6t $T=4816 942 0 0 $X=4792 $Y=942
XX246034E0159 GND! VDD! GND! BLB<8> 115 296 BL<8> WL<0> 295 114 297 
+	WL<1> 268 268 270 sram_6t $T=4816 18 0 0 $X=4792 $Y=18
XX246034E0160 GND! VDD! GND! BLB<9> 139 305 BL<9> WL<0> 304 138 306 
+	WL<1> 268 268 270 sram_6t $T=5320 18 0 0 $X=5296 $Y=18
XX246034E0161 GND! VDD! GND! BLB<11> 137 308 BL<11> WL<0> 307 136 309 
+	WL<1> 268 268 270 sram_6t $T=6328 18 0 0 $X=6304 $Y=18
XX246034E0162 GND! VDD! GND! BLB<10> 135 311 BL<10> WL<0> 310 134 312 
+	WL<1> 268 268 270 sram_6t $T=5824 18 0 0 $X=5800 $Y=18
XX246034E0163 GND! VDD! GND! BLB<1> 65 50 BL<1> WL<3> WL<2> 64 51 
+	WL<4> 268 268 272 sram_6t $T=616 2790 0 0 $X=592 $Y=2790
XX246034E0164 GND! VDD! GND! BLB<0> 67 46 BL<0> WL<3> WL<2> 66 47 
+	WL<4> 268 268 272 sram_6t $T=112 2790 0 0 $X=88 $Y=2790
XX246034E0165 GND! VDD! GND! BLB<14> 171 314 BL<14> WL<0> 313 170 315 
+	WL<1> 268 268 270 sram_6t $T=8176 18 0 0 $X=8152 $Y=18
XX246034E0166 GND! VDD! GND! BLB<15> 169 317 BL<15> WL<0> 316 168 318 
+	WL<1> 268 268 270 sram_6t $T=8680 18 0 0 $X=8656 $Y=18
XX246034E0167 GND! VDD! GND! BLB<13> 167 320 BL<13> WL<0> 319 166 321 
+	WL<1> 268 268 270 sram_6t $T=7672 18 0 0 $X=7648 $Y=18
XX246034E0168 GND! VDD! GND! BLB<12> 165 323 BL<12> WL<0> 322 164 324 
+	WL<1> 268 268 270 sram_6t $T=7168 18 0 0 $X=7144 $Y=18
XX246034E0169 GND! VDD! GND! BLB<4> 89 287 BL<4> WL<0> 286 88 288 
+	WL<1> 268 268 270 sram_6t $T=2464 18 0 0 $X=2440 $Y=18
XX246034E0170 GND! VDD! GND! BLB<5> 87 290 BL<5> WL<0> 289 86 291 
+	WL<1> 268 268 270 sram_6t $T=2968 18 0 0 $X=2944 $Y=18
XX246034E0171 GND! VDD! GND! BLB<7> 113 299 BL<7> WL<0> 298 112 300 
+	WL<1> 268 268 270 sram_6t $T=3976 18 0 0 $X=3952 $Y=18
XX246034E0172 GND! VDD! GND! BLB<6> 111 302 BL<6> WL<0> 301 110 303 
+	WL<1> 268 268 270 sram_6t $T=3472 18 0 0 $X=3448 $Y=18
XX246034E0173 GND! VDD! GND! BLB<2> 61 278 BL<2> WL<0> 277 60 279 
+	WL<1> 268 268 270 sram_6t $T=1120 18 0 0 $X=1096 $Y=18
XX246034E0174 GND! VDD! GND! BLB<3> 85 293 BL<3> WL<0> 292 84 294 
+	WL<1> 268 268 270 sram_6t $T=1624 18 0 0 $X=1600 $Y=18
XX246034E0175 GND! VDD! GND! BLB<1> 59 281 BL<1> WL<0> 280 58 282 
+	WL<1> 268 268 270 sram_6t $T=616 18 0 0 $X=592 $Y=18
XX246034E0176 GND! VDD! GND! BLB<0> 57 284 BL<0> WL<0> 283 56 285 
+	WL<1> 268 268 270 sram_6t $T=112 18 0 0 $X=88 $Y=18
.ends memory_array_8by16
