* PEX netlist file	Sat Apr 12 19:00:40 2025	invx4
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 0

* Top of hierarchy  cell=invx4
.subckt invx4 GND! VDD! OUT IN
*.floating_nets 6 7 _GENERATED_8 _GENERATED_9 _GENERATED_10
MM1 GND! IN OUT nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=414 $Y=295  $PIN_XY=444,210,414,295,384,210 $DEVICE_ID=1001
MM2 OUT IN GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=246 $Y=295  $PIN_XY=276,210,246,295,216,210 $DEVICE_ID=1001
MM3 VDD! IN OUT pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=750 $Y=397  $PIN_XY=780,380,750,397,720,380 $DEVICE_ID=1003
MM4 OUT IN VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=582 $Y=397  $PIN_XY=612,380,582,397,552,380 $DEVICE_ID=1003
MM5 VDD! IN OUT pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=414 $Y=295  $PIN_XY=444,380,414,295,384,380 $DEVICE_ID=1003
MM6 OUT IN VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=246 $Y=295  $PIN_XY=276,380,246,295,216,380 $DEVICE_ID=1003
.ends invx4
