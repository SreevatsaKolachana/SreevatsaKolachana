* PEX netlist file	Thu Apr 17 16:10:37 2025	read_circuit
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 1
.subckt inv 2 3 4 5 7 8 9
*.floating_nets 6 10 11 12
MM1 4 5 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=222 $Y=294  $PIN_XY=252,210,222,294,192,210 $DEVICE_ID=1001
MM2 3 5 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=390 $Y=395  $PIN_XY=420,380,390,395,360,380 $DEVICE_ID=1003
MM3 4 5 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=222 $Y=294  $PIN_XY=252,380,222,294,192,380 $DEVICE_ID=1003
.ends inv
.subckt nand 2 3 4 5 6 10 11 12
*.floating_nets 8 9 13 14 15 16
MM1 4 6 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=808 $Y=522  $PIN_XY=838,438,808,522,778,438 $DEVICE_ID=1001
MM2 7 5 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=640 $Y=522  $PIN_XY=670,438,640,522,610,438 $DEVICE_ID=1001
MM3 3 6 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=808 $Y=522  $PIN_XY=838,608,808,522,778,608 $DEVICE_ID=1003
MM4 4 5 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=640 $Y=522  $PIN_XY=670,608,640,522,610,608 $DEVICE_ID=1003
.ends nand
.subckt invx4 2 3 4 5 6 7 8
*.floating_nets 9 10 11 12 13 14 15 16 17 18
MM1 2 5 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=414 $Y=294  $PIN_XY=444,210,414,294,384,210 $DEVICE_ID=1001
MM2 4 5 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=246 $Y=294  $PIN_XY=276,210,246,294,216,210 $DEVICE_ID=1001
MM3 3 5 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=750 $Y=395  $PIN_XY=780,380,750,395,720,380 $DEVICE_ID=1003
MM4 4 5 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=582 $Y=395  $PIN_XY=612,380,582,395,552,380 $DEVICE_ID=1003
MM5 3 5 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=414 $Y=294  $PIN_XY=444,380,414,294,384,380 $DEVICE_ID=1003
MM6 4 5 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=246 $Y=294  $PIN_XY=276,380,246,294,216,380 $DEVICE_ID=1003
.ends invx4

* Hierarchy Level 0

* Top of hierarchy  cell=read_circuit
.subckt read_circuit BLBAR 5 BL 7 OUT
XXE1FF984B1 2 3 5 BLBAR 9 10 11 invx4 $T=-24 4 0 0 $X=0 $Y=4
XXE1FF984B2 2 3 7 5 BL 9 10 11 nand $T=422 -224 0 0 $X=840 $Y=4
XXE1FF984B3 2 3 OUT 7 9 10 11 inv $T=1512 4 0 0 $X=1512 $Y=4
.ends read_circuit
