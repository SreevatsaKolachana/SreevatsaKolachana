package i2cmb_env_pkg;
    import ncsu_pkg::*;
    import data_pkg::*;
    import i2c_pkg::*;
    import wb_pkg::*;
    `include "../../ncsu_pkg/ncsu_macros.svh"
    `include "src/i2cmb_env_configuration.svh"
    `include "src/i2cmb_coverage.svh"
    `include "src/i2cmb_scoreboard.svh"
    `include "src/i2cmb_predictor.svh"
    `include "src/i2cmb_generator.svh"
    `include "src/i2cmb_environment.svh"
    `include "src/i2cmb_test.svh"
    `include "src/test_i2cmb_reg_addrs.svh"
    `include "src/test_i2cmb_reg_defaults.svh"
    `include "src/test_i2cmb_reg_faultaddrs.svh"
    `include "src/test_i2cmb_reg_transactions.svh"
    `include "src/test_i2cmb_reg_writeouts.svh"
    `include "src/test_i2cmbFSM_before.svh"
    `include "src/test_i2cmbFSM_starts.svh"
    `include "src/test_i2cmbFSM_stops.svh"
    `include "src/test_i2cmbFSM_writefirst.svh"
    `include "src/test_i2cmbFSM_bus_ranges.svh"
    `include "src/test_i2cmb_random.svh"
endpackage