* PEX netlist file	Tue Apr 15 19:44:05 2025	nand
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 0

* Top of hierarchy  cell=nand
.subckt nand GND! VDD! Y A B 7 8 9
*.floating_nets 10 11 12 13 _GENERATED_14 _GENERATED_15 _GENERATED_16
MM1 Y B 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=808 $Y=522  $PIN_XY=838,438,808,522,778,438 $DEVICE_ID=1001
MM2 7 A GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=640 $Y=522  $PIN_XY=670,438,640,522,610,438 $DEVICE_ID=1001
MM3 VDD! B Y pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=808 $Y=522  $PIN_XY=838,608,808,522,778,608 $DEVICE_ID=1003
MM4 Y A VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=640 $Y=522  $PIN_XY=670,608,640,522,610,608 $DEVICE_ID=1003
.ends nand
