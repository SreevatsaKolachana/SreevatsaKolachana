* PEX netlist file	Thu Apr 17 14:29:52 2025	nor
* icv_netlist Version RHEL64 W-2024.09-SP2.11100136 2024/12/03
*.UNIT=4000

* Hierarchy Level 0

* Top of hierarchy  cell=nor
.subckt nor GND! VDD! Y A B 7
*.floating_nets 8 9 10 11 _GENERATED_12 _GENERATED_13 _GENERATED_14
MM1 GND! B Y nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1018 $Y=296  $PIN_XY=1048,212,1018,296,988,212 $DEVICE_ID=1001
MM2 Y A GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=850 $Y=296  $PIN_XY=880,212,850,296,820,212 $DEVICE_ID=1001
MM3 Y B 7 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1018 $Y=296  $PIN_XY=1048,382,1018,296,988,382 $DEVICE_ID=1003
MM4 7 A VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=850 $Y=296  $PIN_XY=880,382,850,296,820,382 $DEVICE_ID=1003
.ends nor
